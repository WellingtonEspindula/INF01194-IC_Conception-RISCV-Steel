
module iopads(clock, reset, halt, 
	rw_address,
	read_data,
	read_request,
	read_response,
	write_data,
	write_strobe,
	write_request,
	write_response,
	irq_external,
	irq_external_response,
	irq_timer,
	irq_timer_response,
	irq_software,
	irq_software_response,
	irq_fast,
	irq_fast_response,
	real_time_clock,
     rw_address_O,
     clock_I, reset_I, halt_I,
     read_data_I,
     read_request_O,
     read_response_I,
     write_data_O,
     write_strobe_O,
     write_request_O,
     write_response_I,
     irq_external_I,
     irq_external_response_O,
     irq_timer_I,
     irq_timer_response_O,
     irq_software_I,
     irq_software_response_O,
     irq_fast_I,
     irq_fast_response_O,
     real_time_clock_I);

     input clock, reset, halt;
	output [31:0] rw_address;
	input [31:0] read_data;
	output read_request;
	input read_response;
	output [31:0] write_data;
	output [3:0] write_strobe;
	output write_request;
     input write_response;
     input irq_external;
	output irq_external_response;
	input irq_timer;
	output irq_timer_response;
	input irq_software;
	output irq_software_response;
	input [15:0] irq_fast;
	output [15:0] irq_fast_response;
     input  [63:0] real_time_clock;

     output clock_I, reset_I, halt_I;
     input [31:0]  rw_address_O;
     output  [31:0]  read_data_I;
     input read_request_O;
     output  read_response_I;
     input [31:0]  write_data_O;
     input [3:0 ]  write_strobe_O;
     input write_request_O;
     output  write_response_I;
     output  irq_external_I;
     input irq_external_response_O;
     output  irq_timer_I;
     input irq_timer_response_O;
     output  irq_software_I;
     input irq_software_response_O;
     output  [15:0]  irq_fast_I;
     input [15:0]  irq_fast_response_O;
     output  [63:0]  real_time_clock_I;

     ICP PAD_clk_i(.PAD(clock), .Y(clock_I));
     ICP PAD_reset_i(.PAD(reset), .Y(reset_I));
     ICP PAD_halt_i(.PAD(halt), .Y(halt_I));

     BD8P PAD_rw_address_o_0(.A(rw_address_O[0]), .PAD(rw_address[0]));
     BD8P PAD_rw_address_o_1(.A(rw_address_O[1]), .PAD(rw_address[1]));
     BD8P PAD_rw_address_o_2(.A(rw_address_O[2]), .PAD(rw_address[2]));
     BD8P PAD_rw_address_o_3(.A(rw_address_O[3]), .PAD(rw_address[3]));
     BD8P PAD_rw_address_o_4(.A(rw_address_O[4]), .PAD(rw_address[4]));
     BD8P PAD_rw_address_o_5(.A(rw_address_O[5]), .PAD(rw_address[5]));
     BD8P PAD_rw_address_o_6(.A(rw_address_O[6]), .PAD(rw_address[6]));
     BD8P PAD_rw_address_o_7(.A(rw_address_O[7]), .PAD(rw_address[7]));
     BD8P PAD_rw_address_o_8(.A(rw_address_O[8]), .PAD(rw_address[8]));
     BD8P PAD_rw_address_o_9(.A(rw_address_O[9]), .PAD(rw_address[9]));
     BD8P PAD_rw_address_o_10(.A(rw_address_O[10]), .PAD(rw_address[10]));
     BD8P PAD_rw_address_o_11(.A(rw_address_O[11]), .PAD(rw_address[11]));
     BD8P PAD_rw_address_o_12(.A(rw_address_O[12]), .PAD(rw_address[12]));
     BD8P PAD_rw_address_o_13(.A(rw_address_O[13]), .PAD(rw_address[13]));
     BD8P PAD_rw_address_o_14(.A(rw_address_O[14]), .PAD(rw_address[14]));
     BD8P PAD_rw_address_o_15(.A(rw_address_O[15]), .PAD(rw_address[15]));
     BD8P PAD_rw_address_o_16(.A(rw_address_O[16]), .PAD(rw_address[16]));
     BD8P PAD_rw_address_o_17(.A(rw_address_O[17]), .PAD(rw_address[17]));
     BD8P PAD_rw_address_o_18(.A(rw_address_O[18]), .PAD(rw_address[18]));
     BD8P PAD_rw_address_o_19(.A(rw_address_O[19]), .PAD(rw_address[19]));
     BD8P PAD_rw_address_o_20(.A(rw_address_O[20]), .PAD(rw_address[20]));
     BD8P PAD_rw_address_o_21(.A(rw_address_O[21]), .PAD(rw_address[21]));
     BD8P PAD_rw_address_o_22(.A(rw_address_O[22]), .PAD(rw_address[22]));
     BD8P PAD_rw_address_o_23(.A(rw_address_O[23]), .PAD(rw_address[23]));
     BD8P PAD_rw_address_o_24(.A(rw_address_O[24]), .PAD(rw_address[24]));
     BD8P PAD_rw_address_o_25(.A(rw_address_O[25]), .PAD(rw_address[25]));
     BD8P PAD_rw_address_o_26(.A(rw_address_O[26]), .PAD(rw_address[26]));
     BD8P PAD_rw_address_o_27(.A(rw_address_O[27]), .PAD(rw_address[27]));
     BD8P PAD_rw_address_o_28(.A(rw_address_O[28]), .PAD(rw_address[28]));
     BD8P PAD_rw_address_o_29(.A(rw_address_O[29]), .PAD(rw_address[29]));
     BD8P PAD_rw_address_o_30(.A(rw_address_O[30]), .PAD(rw_address[30]));
     BD8P PAD_rw_address_o_31(.A(rw_address_O[31]), .PAD(rw_address[31]));

     ICP PAD_read_data_i_0(.PAD(read_data[0]), .Y(read_data_I[0]));
     ICP PAD_read_data_i_1(.PAD(read_data[1]), .Y(read_data_I[1]));
     ICP PAD_read_data_i_2(.PAD(read_data[2]), .Y(read_data_I[2]));
     ICP PAD_read_data_i_3(.PAD(read_data[3]), .Y(read_data_I[3]));
     ICP PAD_read_data_i_4(.PAD(read_data[4]), .Y(read_data_I[4]));
     ICP PAD_read_data_i_5(.PAD(read_data[5]), .Y(read_data_I[5]));
     ICP PAD_read_data_i_6(.PAD(read_data[6]), .Y(read_data_I[6]));
     ICP PAD_read_data_i_7(.PAD(read_data[7]), .Y(read_data_I[7]));
     ICP PAD_read_data_i_8(.PAD(read_data[8]), .Y(read_data_I[8]));
     ICP PAD_read_data_i_9(.PAD(read_data[9]), .Y(read_data_I[9]));
     ICP PAD_read_data_i_10(.PAD(read_data[10]), .Y(read_data_I[10]));
     ICP PAD_read_data_i_11(.PAD(read_data[11]), .Y(read_data_I[11]));
     ICP PAD_read_data_i_12(.PAD(read_data[12]), .Y(read_data_I[12]));
     ICP PAD_read_data_i_13(.PAD(read_data[13]), .Y(read_data_I[13]));
     ICP PAD_read_data_i_14(.PAD(read_data[14]), .Y(read_data_I[14]));
     ICP PAD_read_data_i_15(.PAD(read_data[15]), .Y(read_data_I[15]));
     ICP PAD_read_data_i_16(.PAD(read_data[16]), .Y(read_data_I[16]));
     ICP PAD_read_data_i_17(.PAD(read_data[17]), .Y(read_data_I[17]));
     ICP PAD_read_data_i_18(.PAD(read_data[18]), .Y(read_data_I[18]));
     ICP PAD_read_data_i_19(.PAD(read_data[19]), .Y(read_data_I[19]));
     ICP PAD_read_data_i_20(.PAD(read_data[20]), .Y(read_data_I[20]));
     ICP PAD_read_data_i_21(.PAD(read_data[21]), .Y(read_data_I[21]));
     ICP PAD_read_data_i_22(.PAD(read_data[22]), .Y(read_data_I[22]));
     ICP PAD_read_data_i_23(.PAD(read_data[23]), .Y(read_data_I[23]));
     ICP PAD_read_data_i_24(.PAD(read_data[24]), .Y(read_data_I[24]));
     ICP PAD_read_data_i_25(.PAD(read_data[25]), .Y(read_data_I[25]));
     ICP PAD_read_data_i_26(.PAD(read_data[26]), .Y(read_data_I[26]));
     ICP PAD_read_data_i_27(.PAD(read_data[27]), .Y(read_data_I[27]));
     ICP PAD_read_data_i_28(.PAD(read_data[28]), .Y(read_data_I[28]));
     ICP PAD_read_data_i_29(.PAD(read_data[29]), .Y(read_data_I[29]));
     ICP PAD_read_data_i_30(.PAD(read_data[30]), .Y(read_data_I[30]));
     ICP PAD_read_data_i_31(.PAD(read_data[31]), .Y(read_data_I[31]));

     BD8P PAD_read_request_o(.A(read_request_O), .PAD(read_request));
     ICP PAD_read_response_i(.PAD(read_response), .Y(read_response_I));

     BD8P PAD_write_data_o_0(.A(write_data_O[0]), .PAD(write_data[0]));
     BD8P PAD_write_data_o_1(.A(write_data_O[1]), .PAD(write_data[1]));
     BD8P PAD_write_data_o_2(.A(write_data_O[2]), .PAD(write_data[2]));
     BD8P PAD_write_data_o_3(.A(write_data_O[3]), .PAD(write_data[3]));
     BD8P PAD_write_data_o_4(.A(write_data_O[4]), .PAD(write_data[4]));
     BD8P PAD_write_data_o_5(.A(write_data_O[5]), .PAD(write_data[5]));
     BD8P PAD_write_data_o_6(.A(write_data_O[6]), .PAD(write_data[6]));
     BD8P PAD_write_data_o_7(.A(write_data_O[7]), .PAD(write_data[7]));
     BD8P PAD_write_data_o_8(.A(write_data_O[8]), .PAD(write_data[8]));
     BD8P PAD_write_data_o_9(.A(write_data_O[9]), .PAD(write_data[9]));
     BD8P PAD_write_data_o_10(.A(write_data_O[10]), .PAD(write_data[10]));
     BD8P PAD_write_data_o_11(.A(write_data_O[11]), .PAD(write_data[11]));
     BD8P PAD_write_data_o_12(.A(write_data_O[12]), .PAD(write_data[12]));
     BD8P PAD_write_data_o_13(.A(write_data_O[13]), .PAD(write_data[13]));
     BD8P PAD_write_data_o_14(.A(write_data_O[14]), .PAD(write_data[14]));
     BD8P PAD_write_data_o_15(.A(write_data_O[15]), .PAD(write_data[15]));
     BD8P PAD_write_data_o_16(.A(write_data_O[16]), .PAD(write_data[16]));
     BD8P PAD_write_data_o_17(.A(write_data_O[17]), .PAD(write_data[17]));
     BD8P PAD_write_data_o_18(.A(write_data_O[18]), .PAD(write_data[18]));
     BD8P PAD_write_data_o_19(.A(write_data_O[19]), .PAD(write_data[19]));
     BD8P PAD_write_data_o_20(.A(write_data_O[20]), .PAD(write_data[20]));
     BD8P PAD_write_data_o_21(.A(write_data_O[21]), .PAD(write_data[21]));
     BD8P PAD_write_data_o_22(.A(write_data_O[22]), .PAD(write_data[22]));
     BD8P PAD_write_data_o_23(.A(write_data_O[23]), .PAD(write_data[23]));
     BD8P PAD_write_data_o_24(.A(write_data_O[24]), .PAD(write_data[24]));
     BD8P PAD_write_data_o_25(.A(write_data_O[25]), .PAD(write_data[25]));
     BD8P PAD_write_data_o_26(.A(write_data_O[26]), .PAD(write_data[26]));
     BD8P PAD_write_data_o_27(.A(write_data_O[27]), .PAD(write_data[27]));
     BD8P PAD_write_data_o_28(.A(write_data_O[28]), .PAD(write_data[28]));
     BD8P PAD_write_data_o_29(.A(write_data_O[29]), .PAD(write_data[29]));
     BD8P PAD_write_data_o_30(.A(write_data_O[30]), .PAD(write_data[30]));
     BD8P PAD_write_data_o_31(.A(write_data_O[31]), .PAD(write_data[31]));

     BD8P PAD_write_strobe_o_0(.A(write_strobe_O[0]), .PAD(write_strobe[0]));
     BD8P PAD_write_strobe_o_1(.A(write_strobe_O[1]), .PAD(write_strobe[1]));
     BD8P PAD_write_strobe_o_2(.A(write_strobe_O[2]), .PAD(write_strobe[2]));
     BD8P PAD_write_strobe_o_3(.A(write_strobe_O[3]), .PAD(write_strobe[3]));
     
     BD8P PAD_write_request_o(.A(write_request_O), .PAD(write_request));
     ICP PAD_write_response_i(.PAD(write_response), .Y(write_response_I));

     ICP PAD_irq_external_i(.PAD(irq_external), .Y(irq_external_I));
     BD8P PAD_irq_external_response_o(.A(irq_external_response_O), .PAD(irq_external_response));

     ICP PAD_irq_timer_i(.PAD(irq_timer), .Y(irq_timer_I));
     BD8P PAD_irq_timer_response_o(.A(irq_timer_response_O), .PAD(irq_timer_response));

     ICP PAD_irq_software_i(.PAD(irq_software), .Y(irq_software_I));
     BD8P PAD_irq_software_response_o(.A(irq_software_response_O), .PAD(irq_software_response));
     
     ICP PAD_irq_fast_i_0(.PAD(irq_fast[0]), .Y(irq_fast_I[0]));
     ICP PAD_irq_fast_i_1(.PAD(irq_fast[1]), .Y(irq_fast_I[1]));
     ICP PAD_irq_fast_i_2(.PAD(irq_fast[2]), .Y(irq_fast_I[2]));
     ICP PAD_irq_fast_i_3(.PAD(irq_fast[3]), .Y(irq_fast_I[3]));
     ICP PAD_irq_fast_i_4(.PAD(irq_fast[4]), .Y(irq_fast_I[4]));
     ICP PAD_irq_fast_i_5(.PAD(irq_fast[5]), .Y(irq_fast_I[5]));
     ICP PAD_irq_fast_i_6(.PAD(irq_fast[6]), .Y(irq_fast_I[6]));
     ICP PAD_irq_fast_i_7(.PAD(irq_fast[7]), .Y(irq_fast_I[7]));
     ICP PAD_irq_fast_i_8(.PAD(irq_fast[8]), .Y(irq_fast_I[8]));
     ICP PAD_irq_fast_i_9(.PAD(irq_fast[9]), .Y(irq_fast_I[9]));
     ICP PAD_irq_fast_i_10(.PAD(irq_fast[10]), .Y(irq_fast_I[10]));
     ICP PAD_irq_fast_i_11(.PAD(irq_fast[11]), .Y(irq_fast_I[11]));
     ICP PAD_irq_fast_i_12(.PAD(irq_fast[12]), .Y(irq_fast_I[12]));
     ICP PAD_irq_fast_i_13(.PAD(irq_fast[13]), .Y(irq_fast_I[13]));
     ICP PAD_irq_fast_i_14(.PAD(irq_fast[14]), .Y(irq_fast_I[14]));
     ICP PAD_irq_fast_i_15(.PAD(irq_fast[15]), .Y(irq_fast_I[15]));

     BD8P PAD_irq_fast_response_o_0(.A(irq_fast_response_O[0]), .PAD(irq_fast_response[0]));
     BD8P PAD_irq_fast_response_o_1(.A(irq_fast_response_O[1]), .PAD(irq_fast_response[1]));
     BD8P PAD_irq_fast_response_o_2(.A(irq_fast_response_O[2]), .PAD(irq_fast_response[2]));
     BD8P PAD_irq_fast_response_o_3(.A(irq_fast_response_O[3]), .PAD(irq_fast_response[3]));
     BD8P PAD_irq_fast_response_o_4(.A(irq_fast_response_O[4]), .PAD(irq_fast_response[4]));
     BD8P PAD_irq_fast_response_o_5(.A(irq_fast_response_O[5]), .PAD(irq_fast_response[5]));
     BD8P PAD_irq_fast_response_o_6(.A(irq_fast_response_O[6]), .PAD(irq_fast_response[6]));
     BD8P PAD_irq_fast_response_o_7(.A(irq_fast_response_O[7]), .PAD(irq_fast_response[7]));
     BD8P PAD_irq_fast_response_o_8(.A(irq_fast_response_O[8]), .PAD(irq_fast_response[8]));
     BD8P PAD_irq_fast_response_o_9(.A(irq_fast_response_O[9]), .PAD(irq_fast_response[9]));
     BD8P PAD_irq_fast_response_o_10(.A(irq_fast_response_O[10]), .PAD(irq_fast_response[10]));
     BD8P PAD_irq_fast_response_o_11(.A(irq_fast_response_O[11]), .PAD(irq_fast_response[11]));
     BD8P PAD_irq_fast_response_o_12(.A(irq_fast_response_O[12]), .PAD(irq_fast_response[12]));
     BD8P PAD_irq_fast_response_o_13(.A(irq_fast_response_O[13]), .PAD(irq_fast_response[13]));
     BD8P PAD_irq_fast_response_o_14(.A(irq_fast_response_O[14]), .PAD(irq_fast_response[14]));
     BD8P PAD_irq_fast_response_o_15(.A(irq_fast_response_O[15]), .PAD(irq_fast_response[15]));

     ICP PAD_real_time_clock_i_0(.PAD(real_time_clock[0]), .Y(real_time_clock_I[0]));
     ICP PAD_real_time_clock_i_1(.PAD(real_time_clock[1]), .Y(real_time_clock_I[1]));
     ICP PAD_real_time_clock_i_2(.PAD(real_time_clock[2]), .Y(real_time_clock_I[2]));
     ICP PAD_real_time_clock_i_3(.PAD(real_time_clock[3]), .Y(real_time_clock_I[3]));
     ICP PAD_real_time_clock_i_4(.PAD(real_time_clock[4]), .Y(real_time_clock_I[4]));
     ICP PAD_real_time_clock_i_5(.PAD(real_time_clock[5]), .Y(real_time_clock_I[5]));
     ICP PAD_real_time_clock_i_6(.PAD(real_time_clock[6]), .Y(real_time_clock_I[6]));
     ICP PAD_real_time_clock_i_7(.PAD(real_time_clock[7]), .Y(real_time_clock_I[7]));
     ICP PAD_real_time_clock_i_8(.PAD(real_time_clock[8]), .Y(real_time_clock_I[8]));
     ICP PAD_real_time_clock_i_9(.PAD(real_time_clock[9]), .Y(real_time_clock_I[9]));
     ICP PAD_real_time_clock_i_10(.PAD(real_time_clock[10]), .Y(real_time_clock_I[10]));
     ICP PAD_real_time_clock_i_11(.PAD(real_time_clock[11]), .Y(real_time_clock_I[11]));
     ICP PAD_real_time_clock_i_12(.PAD(real_time_clock[12]), .Y(real_time_clock_I[12]));
     ICP PAD_real_time_clock_i_13(.PAD(real_time_clock[13]), .Y(real_time_clock_I[13]));
     ICP PAD_real_time_clock_i_14(.PAD(real_time_clock[14]), .Y(real_time_clock_I[14]));
     ICP PAD_real_time_clock_i_15(.PAD(real_time_clock[15]), .Y(real_time_clock_I[15]));
     ICP PAD_real_time_clock_i_16(.PAD(real_time_clock[16]), .Y(real_time_clock_I[16]));
     ICP PAD_real_time_clock_i_17(.PAD(real_time_clock[17]), .Y(real_time_clock_I[17]));
     ICP PAD_real_time_clock_i_18(.PAD(real_time_clock[18]), .Y(real_time_clock_I[18]));
     ICP PAD_real_time_clock_i_19(.PAD(real_time_clock[19]), .Y(real_time_clock_I[19]));
     ICP PAD_real_time_clock_i_20(.PAD(real_time_clock[20]), .Y(real_time_clock_I[20]));
     ICP PAD_real_time_clock_i_21(.PAD(real_time_clock[21]), .Y(real_time_clock_I[21]));
     ICP PAD_real_time_clock_i_22(.PAD(real_time_clock[22]), .Y(real_time_clock_I[22]));
     ICP PAD_real_time_clock_i_23(.PAD(real_time_clock[23]), .Y(real_time_clock_I[23]));
     ICP PAD_real_time_clock_i_24(.PAD(real_time_clock[24]), .Y(real_time_clock_I[24]));
     ICP PAD_real_time_clock_i_25(.PAD(real_time_clock[25]), .Y(real_time_clock_I[25]));
     ICP PAD_real_time_clock_i_26(.PAD(real_time_clock[26]), .Y(real_time_clock_I[26]));
     ICP PAD_real_time_clock_i_27(.PAD(real_time_clock[27]), .Y(real_time_clock_I[27]));
     ICP PAD_real_time_clock_i_28(.PAD(real_time_clock[28]), .Y(real_time_clock_I[28]));
     ICP PAD_real_time_clock_i_29(.PAD(real_time_clock[29]), .Y(real_time_clock_I[29]));
     ICP PAD_real_time_clock_i_30(.PAD(real_time_clock[30]), .Y(real_time_clock_I[30]));
     ICP PAD_real_time_clock_i_31(.PAD(real_time_clock[31]), .Y(real_time_clock_I[31]));
     ICP PAD_real_time_clock_i_32(.PAD(real_time_clock[32]), .Y(real_time_clock_I[32]));
     ICP PAD_real_time_clock_i_33(.PAD(real_time_clock[33]), .Y(real_time_clock_I[33]));
     ICP PAD_real_time_clock_i_34(.PAD(real_time_clock[34]), .Y(real_time_clock_I[34]));
     ICP PAD_real_time_clock_i_35(.PAD(real_time_clock[35]), .Y(real_time_clock_I[35]));
     ICP PAD_real_time_clock_i_36(.PAD(real_time_clock[36]), .Y(real_time_clock_I[36]));
     ICP PAD_real_time_clock_i_37(.PAD(real_time_clock[37]), .Y(real_time_clock_I[37]));
     ICP PAD_real_time_clock_i_38(.PAD(real_time_clock[38]), .Y(real_time_clock_I[38]));
     ICP PAD_real_time_clock_i_39(.PAD(real_time_clock[39]), .Y(real_time_clock_I[39]));
     ICP PAD_real_time_clock_i_40(.PAD(real_time_clock[40]), .Y(real_time_clock_I[40]));
     ICP PAD_real_time_clock_i_41(.PAD(real_time_clock[41]), .Y(real_time_clock_I[41]));
     ICP PAD_real_time_clock_i_42(.PAD(real_time_clock[42]), .Y(real_time_clock_I[42]));
     ICP PAD_real_time_clock_i_43(.PAD(real_time_clock[43]), .Y(real_time_clock_I[43]));
     ICP PAD_real_time_clock_i_44(.PAD(real_time_clock[44]), .Y(real_time_clock_I[44]));
     ICP PAD_real_time_clock_i_45(.PAD(real_time_clock[45]), .Y(real_time_clock_I[45]));
     ICP PAD_real_time_clock_i_46(.PAD(real_time_clock[46]), .Y(real_time_clock_I[46]));
     ICP PAD_real_time_clock_i_47(.PAD(real_time_clock[47]), .Y(real_time_clock_I[47]));
     ICP PAD_real_time_clock_i_48(.PAD(real_time_clock[48]), .Y(real_time_clock_I[48]));
     ICP PAD_real_time_clock_i_49(.PAD(real_time_clock[49]), .Y(real_time_clock_I[49]));
     ICP PAD_real_time_clock_i_50(.PAD(real_time_clock[50]), .Y(real_time_clock_I[50]));
     ICP PAD_real_time_clock_i_51(.PAD(real_time_clock[51]), .Y(real_time_clock_I[51]));
     ICP PAD_real_time_clock_i_52(.PAD(real_time_clock[52]), .Y(real_time_clock_I[52]));
     ICP PAD_real_time_clock_i_53(.PAD(real_time_clock[53]), .Y(real_time_clock_I[53]));
     ICP PAD_real_time_clock_i_54(.PAD(real_time_clock[54]), .Y(real_time_clock_I[54]));
     ICP PAD_real_time_clock_i_55(.PAD(real_time_clock[55]), .Y(real_time_clock_I[55]));
     ICP PAD_real_time_clock_i_56(.PAD(real_time_clock[56]), .Y(real_time_clock_I[56]));
     ICP PAD_real_time_clock_i_57(.PAD(real_time_clock[57]), .Y(real_time_clock_I[57]));
     ICP PAD_real_time_clock_i_58(.PAD(real_time_clock[58]), .Y(real_time_clock_I[58]));
     ICP PAD_real_time_clock_i_59(.PAD(real_time_clock[59]), .Y(real_time_clock_I[59]));
     ICP PAD_real_time_clock_i_60(.PAD(real_time_clock[60]), .Y(real_time_clock_I[60]));
     ICP PAD_real_time_clock_i_61(.PAD(real_time_clock[61]), .Y(real_time_clock_I[61]));
     ICP PAD_real_time_clock_i_62(.PAD(real_time_clock[62]), .Y(real_time_clock_I[62]));
     ICP PAD_real_time_clock_i_63(.PAD(real_time_clock[63]), .Y(real_time_clock_I[63]));

	VDDORPADP PAD_vdd_E();
	VDDPADP PAD_vdd_core_E();

	VDDPADP PAD_vdd_core_N();
	GNDORPADP PAD_vss_core_N();

	GNDORPADP PAD_vss_W();

	GNDORPADP PAD_vss_S();

	CORNERP PAD_corner_ll();
	CORNERP PAD_corner_lr();
	CORNERP PAD_corner_ul();
	CORNERP PAD_corner_ur();	
endmodule

module top(clock, 
              reset, 
              halt, 
              rw_address,
              read_data,
              read_request,
              read_response,
              write_data,
              write_strobe,
              write_request,
              write_response,
              irq_external,
              irq_external_response,
              irq_timer,
              irq_timer_response,
              irq_software,
              irq_software_response,
              irq_fast,
              irq_fast_response,
              real_time_clock);

     input  clock;
     input  reset;
     input  halt;

     output [31:0]  rw_address;
     input [31:0]  read_data;
     output  read_request;
     input  read_response;
     output [31:0]  write_data;
     output [3:0 ]  write_strobe;
     output  write_request;
     input  write_response;

     input  irq_external;
     output  irq_external_response;
     input  irq_timer;
     output  irq_timer_response;
     input  irq_software;
     output  irq_software_response;
     input [15:0]  irq_fast;
     output [15:0]  irq_fast_response;

     input [63:0]  real_time_clock;


	wire clock_I, reset_I, halt_I;
	
	wire [31:0]  rw_address_O;
	wire  [31:0]  read_data_I;
	wire read_request_O;
	wire  read_response_I;
	wire [31:0]  write_data_O;
	wire [3:0 ]  write_strobe_O;
	wire write_request_O;

	wire  write_response_I;

	wire  irq_external_I;
	wire irq_external_response_O;
	wire  irq_timer_I;
	wire irq_timer_response_O;
	wire  irq_software_I;
	wire irq_software_response_O;
	wire  [15:0]  irq_fast_I;
	wire [15:0]  irq_fast_response_O;

	wire  [63:0]  real_time_clock_I;

	rvsteel_core top_INST(
          .clock(clock_I),
  	     .reset(reset_I),
          .halt(halt_I),
          .rw_address(rw_address_O),
          .read_data(read_data_I),
          .read_request(read_request_O),
          .read_response(read_response_I),
          .write_data(write_data_O),
          .write_strobe(write_strobe_O),
          .write_request(write_request_O),
          .write_response(write_response_I),
          .irq_external(irq_external_I),
          .irq_external_response(irq_external_response_O),
          .irq_timer(irq_timer_I),
          .irq_timer_response(irq_timer_response_O),
          .irq_software(irq_software_I),
          .irq_software_response(irq_software_response_O),
          .irq_fast(irq_fast_I),
          .irq_fast_response(irq_fast_response_O),
          .real_time_clock(real_time_clock_I)
	);

	iopads IOPADS_INST(
          .clock(clock),
          .reset(reset),
          .halt(halt),
          .rw_address(rw_address),
          .read_data(read_data),
          .read_request(read_request),
          .read_response(read_response),
          .write_data(write_data),
          .write_strobe(write_strobe),
          .write_request(write_request),
          .write_response(write_response),
          .irq_external(irq_external),
          .irq_external_response(irq_external_response),
          .irq_timer(irq_timer),
          .irq_timer_response(irq_timer_response),
          .irq_software(irq_software),
          .irq_software_response(irq_software_response),
          .irq_fast(irq_fast),
          .irq_fast_response(irq_fast_response),
          .real_time_clock(real_time_clock),

          .clock_I(clock_I),
          .reset_I(reset_I),
          .halt_I(halt_I),
          .rw_address_O(rw_address_O),
          .read_data_I(read_data_I),
          .read_request_O(read_request_O),
          .read_response_I(read_response_I),
          .write_data_O(write_data_O),
          .write_strobe_O(write_strobe_O),
          .write_request_O(write_request_O),
          .write_response_I(write_response_I),
          .irq_external_I(irq_external_I),
          .irq_external_response_O(irq_external_response_O),
          .irq_timer_I(irq_timer_I),
          .irq_timer_response_O(irq_timer_response_O),
          .irq_software_I(irq_software_I),
          .irq_software_response_O(irq_software_response_O),
          .irq_fast_I(irq_fast_I),
          .irq_fast_response_O(irq_fast_response_O),
          .real_time_clock_I(real_time_clock_I)
	);
endmodule



// Generated by Cadence Genus(TM) Synthesis Solution GENUS15.22 - 15.20-s024_1
// Generated on: Dec 17 2024 07:34:07

// Verification Directory fv/rvsteel_core 

module RC_CG_MOD_AUTO_rvsteel_core(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_9(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_10(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_11(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_12(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_13(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_14(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_15(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_16(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_17(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_18(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_1(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_19(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_20(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_21(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_22(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_23(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_24(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_25(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_26(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_27(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_28(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_2(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_29(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_30(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_31(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_32(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_33(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_34(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_35(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_36(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_37(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_38(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_3(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_39(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_40(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_41(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_4(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_5(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_6(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_7(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_8(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module csa_tree_add_1660_20_group_293(in_0, in_1, in_2, out_0);
  input [31:0] in_0;
  input [33:0] in_1, in_2;
  output [31:0] out_0;
  wire [31:0] in_0;
  wire [33:0] in_1, in_2;
  wire [31:0] out_0;
  wire UNCONNECTED, n_1, n_2, n_3, n_89, n_90, n_92, n_93;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_117, n_118, n_119, n_120;
  wire n_122, n_123, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_147, n_148, n_149;
  wire n_150, n_151, n_152, n_153, n_161, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_246, n_247, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_272, n_273, n_274, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_310, n_311, n_312;
  HAX1 g251(.A (in_1[14]), .B (in_0[14]), .S (n_102), .CO (n_136));
  HAX1 g252(.A (in_1[24]), .B (in_0[24]), .S (n_113), .CO (n_147));
  HAX1 g253(.A (in_1[25]), .B (in_0[25]), .S (n_114), .CO (n_148));
  HAX1 g254(.A (in_1[26]), .B (in_0[26]), .S (n_115), .CO (n_149));
  HAX1 g255(.A (in_1[27]), .B (in_0[27]), .S (n_117), .CO (n_150));
  HAX1 g256(.A (in_1[28]), .B (in_0[28]), .S (n_118), .CO (n_151));
  HAX1 g257(.A (in_1[29]), .B (in_0[29]), .S (n_119), .CO (n_152));
  HAX1 g258(.A (in_1[30]), .B (in_0[30]), .S (n_120), .CO (n_153));
  MU2IX1 g259(.S (in_1[2]), .IN0 (n_2), .IN1 (in_0[2]), .Q (n_89));
  NO2X1 g260(.A (n_3), .B (n_2), .Q (n_122));
  INX1 g261(.A (in_1[2]), .Q (n_3));
  INX1 g262(.A (in_0[2]), .Q (n_2));
  MU2IX1 g263(.S (in_0[3]), .IN0 (n_1), .IN1 (in_1[3]), .Q (n_90));
  NO2I1X1 g264(.B (n_1), .AN (in_0[3]), .Q (n_123));
  INX1 g265(.A (in_1[3]), .Q (n_1));
  HAX1 g266(.A (in_1[15]), .B (in_0[15]), .S (n_103), .CO (n_137));
  HAX2 g270(.A (in_1[5]), .B (in_0[5]), .S (n_92), .CO (n_126));
  HAX1 g271(.A (in_1[6]), .B (in_0[6]), .S (n_93), .CO (n_127));
  HAX1 g272(.A (in_1[7]), .B (in_0[7]), .S (n_95), .CO (n_128));
  HAX1 g273(.A (in_1[8]), .B (in_0[8]), .S (n_96), .CO (n_129));
  HAX1 g274(.A (in_1[9]), .B (in_0[9]), .S (n_97), .CO (n_130));
  HAX1 g275(.A (in_1[10]), .B (in_0[10]), .S (n_98), .CO (n_131));
  HAX1 g276(.A (in_1[11]), .B (in_0[11]), .S (n_99), .CO (n_132));
  HAX1 g277(.A (in_1[12]), .B (in_0[12]), .S (n_100), .CO (n_133));
  HAX1 g278(.A (in_1[13]), .B (in_0[13]), .S (n_101), .CO (n_134));
  HAX1 g279(.A (in_1[16]), .B (in_0[16]), .S (n_104), .CO (n_138));
  HAX1 g280(.A (in_1[17]), .B (in_0[17]), .S (n_106), .CO (n_139));
  HAX1 g281(.A (in_1[18]), .B (in_0[18]), .S (n_107), .CO (n_140));
  HAX1 g282(.A (in_1[19]), .B (in_0[19]), .S (n_108), .CO (n_141));
  HAX1 g283(.A (in_1[20]), .B (in_0[20]), .S (n_109), .CO (n_142));
  HAX1 g284(.A (in_1[21]), .B (in_0[21]), .S (n_110), .CO (n_143));
  HAX1 g285(.A (in_1[22]), .B (in_0[22]), .S (n_111), .CO (n_144));
  HAX1 g286(.A (in_1[23]), .B (in_0[23]), .S (n_112), .CO (n_145));
  NO2X2 g2529(.A (n_300), .B (n_200), .Q (n_301));
  NO2X2 g2531(.A (n_299), .B (n_213), .Q (n_300));
  NO2X4 g2532(.A (n_298), .B (n_196), .Q (n_299));
  NO2X2 g2534(.A (n_297), .B (n_195), .Q (n_298));
  NO2X4 g2535(.A (n_296), .B (n_197), .Q (n_297));
  NO2X4 g2537(.A (n_295), .B (n_198), .Q (n_296));
  NO2X4 g2538(.A (n_294), .B (n_207), .Q (n_295));
  NO2X4 g2540(.A (n_293), .B (n_199), .Q (n_294));
  NO2X4 g2541(.A (n_292), .B (n_201), .Q (n_293));
  NO2X4 g2544(.A (n_304), .B (n_210), .Q (n_292));
  NA2X1 g2547(.A (n_288), .B (n_166), .Q (n_289));
  EN2X1 g2548(.A (n_287), .B (n_223), .Q (out_0[24]));
  NA2X4 g2549(.A (n_287), .B (n_178), .Q (n_288));
  NA2X4 g2550(.A (n_286), .B (n_179), .Q (n_287));
  EN2X1 g2551(.A (n_283), .B (n_216), .Q (out_0[23]));
  NA2X4 g2552(.A (n_285), .B (n_182), .Q (n_286));
  NA2X4 g2553(.A (n_284), .B (n_170), .Q (n_285));
  NA2X4 g2555(.A (n_282), .B (n_172), .Q (n_284));
  AN21X1 g2556(.A (n_279), .B (n_172), .C (n_169), .Q (n_283));
  EO2X1 g2557(.A (n_279), .B (n_220), .Q (out_0[22]));
  NA2X2 g2558(.A (n_281), .B (n_246), .Q (n_282));
  EN2X0 g2559(.A (n_278), .B (n_232), .Q (out_0[19]));
  NA2X2 g2560(.A (n_277), .B (n_164), .Q (n_281));
  NA2I1X1 g2561(.B (n_193), .AN (n_277), .Q (n_280));
  ON21X1 g2562(.A (n_276), .B (n_237), .C (n_246), .Q (n_279));
  EN2X0 g2563(.A (n_276), .B (n_230), .Q (out_0[20]));
  ON21X1 g2564(.A (n_161), .B (n_189), .C (n_192), .Q (n_278));
  EN2X0 g2565(.A (n_161), .B (n_231), .Q (out_0[18]));
  NO2X2 g2566(.A (n_276), .B (n_194), .Q (n_277));
  EN2X0 g2567(.A (n_274), .B (n_219), .Q (out_0[17]));
  NO2X2 g2568(.A (n_307), .B (n_250), .Q (n_276));
  EO2X0 g2571(.A (n_272), .B (n_229), .Q (out_0[16]));
  AN21X1 g2572(.A (n_272), .B (n_167), .C (n_168), .Q (n_274));
  NA2X4 g2573(.A (n_272), .B (n_224), .Q (n_273));
  EO2X0 g2574(.A (n_270), .B (n_234), .Q (out_0[15]));
  NA2X4 g2575(.A (n_271), .B (n_212), .Q (n_272));
  NA2X4 g2576(.A (n_270), .B (n_208), .Q (n_271));
  NA2X4 g2577(.A (n_269), .B (n_211), .Q (n_270));
  EN2X0 g2578(.A (n_268), .B (n_233), .Q (out_0[14]));
  NA2X4 g2579(.A (n_268), .B (n_209), .Q (n_269));
  NA2X4 g2580(.A (n_267), .B (n_186), .Q (n_268));
  EN2X0 g2581(.A (n_266), .B (n_218), .Q (out_0[13]));
  NA2X4 g2582(.A (n_266), .B (n_177), .Q (n_267));
  NA2X4 g2583(.A (n_265), .B (n_181), .Q (n_266));
  EN2X0 g2584(.A (n_264), .B (n_222), .Q (out_0[12]));
  NA2X4 g2585(.A (n_264), .B (n_184), .Q (n_265));
  NA2X4 g2586(.A (n_263), .B (n_203), .Q (n_264));
  EN2X0 g2587(.A (n_262), .B (n_236), .Q (out_0[11]));
  NA2X4 g2588(.A (n_262), .B (n_206), .Q (n_263));
  NA2X4 g2589(.A (n_261), .B (n_202), .Q (n_262));
  EN2X0 g2590(.A (n_260), .B (n_221), .Q (out_0[9]));
  EN2X0 g2591(.A (n_259), .B (n_235), .Q (out_0[10]));
  NA2X4 g2592(.A (n_259), .B (n_205), .Q (n_261));
  AN21X1 g2593(.A (n_257), .B (n_173), .C (n_175), .Q (n_260));
  NA2X2 g2594(.A (n_308), .B (n_247), .Q (n_259));
  EN2X0 g2595(.A (n_257), .B (n_217), .Q (out_0[8]));
  FAX2 g2597(.A (n_127), .B (n_95), .CI (n_256), .S (out_0[7]), .CO
       (n_257));
  FAX2 g2598(.A (n_126), .B (n_93), .CI (n_255), .S (out_0[6]), .CO
       (n_256));
  FAX2 g2599(.A (n_311), .B (n_92), .CI (n_254), .S (out_0[5]), .CO
       (n_255));
  FAX2 g2600(.A (n_123), .B (n_312), .CI (n_253), .S (out_0[4]), .CO
       (n_254));
  FAX2 g2601(.A (n_122), .B (n_90), .CI (n_252), .S (out_0[3]), .CO
       (n_253));
  NO2I1X2 g2603(.B (n_251), .AN (n_89), .Q (n_252));
  OA21X4 g2606(.A (n_306), .B (n_185), .C (n_183), .Q (n_251));
  ON21X1 g2607(.A (n_249), .B (n_191), .C (n_204), .Q (n_250));
  OA21X1 g2609(.A (n_244), .B (n_189), .C (n_192), .Q (n_249));
  AN21X1 g2613(.A (n_174), .B (n_175), .C (n_176), .Q (n_247));
  OA21X1 g2614(.A (n_193), .B (n_165), .C (n_188), .Q (n_246));
  AN21X1 g2617(.A (n_168), .B (n_171), .C (n_180), .Q (n_244));
  OR2X1 g2624(.A (n_194), .B (n_165), .Q (n_237));
  NA2X1 g2625(.A (n_206), .B (n_203), .Q (n_236));
  NA2X1 g2626(.A (n_205), .B (n_202), .Q (n_235));
  AND2X1 g2627(.A (n_208), .B (n_212), .Q (n_234));
  NA2X1 g2628(.A (n_209), .B (n_211), .Q (n_233));
  NO2X1 g2629(.A (n_201), .B (n_210), .Q (n_243));
  NA2I1X1 g2630(.B (n_204), .AN (n_191), .Q (n_232));
  NO2X1 g2631(.A (n_200), .B (n_213), .Q (n_242));
  NO2X1 g2632(.A (n_196), .B (n_195), .Q (n_241));
  NO2X1 g2633(.A (n_197), .B (n_198), .Q (n_240));
  NO2I1X1 g2634(.B (n_189), .AN (n_192), .Q (n_231));
  NO2I1X1 g2635(.B (n_194), .AN (n_193), .Q (n_230));
  NO2X1 g2636(.A (n_207), .B (n_199), .Q (n_239));
  NO2I1X1 g2637(.B (n_168), .AN (n_167), .Q (n_229));
  AND2X1 g2642(.A (n_167), .B (n_171), .Q (n_224));
  NA2X1 g2643(.A (n_164), .B (n_188), .Q (n_228));
  NO2I1X1 g2644(.B (n_190), .AN (n_187), .Q (n_227));
  NA2X1 g2645(.A (n_178), .B (n_166), .Q (n_223));
  NA2X1 g2647(.A (n_184), .B (n_181), .Q (n_222));
  NO2I1X1 g2648(.B (n_176), .AN (n_174), .Q (n_221));
  AND2X1 g2649(.A (n_172), .B (n_170), .Q (n_220));
  NO2I1X1 g2650(.B (n_180), .AN (n_171), .Q (n_219));
  NA2X1 g2651(.A (n_177), .B (n_186), .Q (n_218));
  NA2I1X1 g2652(.B (n_173), .AN (n_175), .Q (n_217));
  AND2X1 g2653(.A (n_182), .B (n_179), .Q (n_216));
  NA2I1X1 g2654(.B (n_183), .AN (n_185), .Q (n_215));
  NO2X1 g2656(.A (n_120), .B (n_152), .Q (n_213));
  NA2X1 g2657(.A (n_103), .B (n_136), .Q (n_212));
  NA2X1 g2658(.A (n_102), .B (n_134), .Q (n_211));
  NO2X1 g2659(.A (n_115), .B (n_148), .Q (n_210));
  OR2X1 g2660(.A (n_102), .B (n_134), .Q (n_209));
  OR2X1 g2661(.A (n_103), .B (n_136), .Q (n_208));
  AND2X1 g2662(.A (n_117), .B (n_149), .Q (n_207));
  OR2X1 g2663(.A (n_99), .B (n_131), .Q (n_206));
  OR2X1 g2664(.A (n_98), .B (n_130), .Q (n_205));
  NA2X1 g2665(.A (n_108), .B (n_140), .Q (n_204));
  NA2X1 g2666(.A (n_99), .B (n_131), .Q (n_203));
  NA2X1 g2667(.A (n_98), .B (n_130), .Q (n_202));
  AND2X1 g2668(.A (n_115), .B (n_148), .Q (n_201));
  AND2X1 g2669(.A (n_120), .B (n_152), .Q (n_200));
  NO2X1 g2670(.A (n_117), .B (n_149), .Q (n_199));
  NO2X1 g2671(.A (n_118), .B (n_150), .Q (n_198));
  AND2X1 g2672(.A (n_118), .B (n_150), .Q (n_197));
  AND2X1 g2673(.A (n_119), .B (n_151), .Q (n_196));
  NO2X1 g2674(.A (n_119), .B (n_151), .Q (n_195));
  NO2X1 g2675(.A (n_109), .B (n_141), .Q (n_194));
  NA2X1 g2676(.A (n_109), .B (n_141), .Q (n_193));
  NA2X1 g2677(.A (n_107), .B (n_139), .Q (n_192));
  NO2X1 g2678(.A (n_108), .B (n_140), .Q (n_191));
  NO2X1 g2679(.A (n_114), .B (n_147), .Q (n_190));
  NO2X1 g2680(.A (n_107), .B (n_139), .Q (n_189));
  INX1 g2681(.A (n_170), .Q (n_169));
  INX1 g2682(.A (n_165), .Q (n_164));
  NA2X1 g2685(.A (n_110), .B (n_142), .Q (n_188));
  NA2X1 g2686(.A (n_114), .B (n_147), .Q (n_187));
  NA2X1 g2687(.A (n_101), .B (n_133), .Q (n_186));
  NO2X1 g2688(.A (in_1[1]), .B (in_0[1]), .Q (n_185));
  OR2X1 g2689(.A (n_100), .B (n_132), .Q (n_184));
  NA2X1 g2690(.A (in_1[1]), .B (in_0[1]), .Q (n_183));
  OR2X1 g2691(.A (n_112), .B (n_144), .Q (n_182));
  NA2X1 g2692(.A (n_132), .B (n_100), .Q (n_181));
  AND2X1 g2693(.A (n_106), .B (n_138), .Q (n_180));
  NA2X1 g2694(.A (n_112), .B (n_144), .Q (n_179));
  OR2X1 g2695(.A (n_113), .B (n_145), .Q (n_178));
  OR2X1 g2696(.A (n_101), .B (n_133), .Q (n_177));
  AND2X1 g2697(.A (n_97), .B (n_129), .Q (n_176));
  AND2X1 g2698(.A (n_96), .B (n_128), .Q (n_175));
  OR2X1 g2699(.A (n_97), .B (n_129), .Q (n_174));
  OR2X1 g2700(.A (n_96), .B (n_128), .Q (n_173));
  OR2X1 g2701(.A (n_111), .B (n_143), .Q (n_172));
  OR2X1 g2702(.A (n_106), .B (n_138), .Q (n_171));
  NA2X1 g2703(.A (n_111), .B (n_143), .Q (n_170));
  AND2X1 g2704(.A (n_137), .B (n_104), .Q (n_168));
  OR2X1 g2705(.A (n_137), .B (n_104), .Q (n_167));
  NA2X1 g2706(.A (n_113), .B (n_145), .Q (n_166));
  NO2X1 g2707(.A (n_110), .B (n_142), .Q (n_165));
  EN2X0 g2(.A (n_251), .B (n_89), .Q (out_0[2]));
  EO2X1 g2709(.A (n_215), .B (n_306), .Q (out_0[1]));
  AND2X1 g2710(.A (n_244), .B (n_273), .Q (n_161));
  EN2X1 g2711(.A (n_304), .B (n_243), .Q (out_0[26]));
  EN2X1 g2712(.A (n_299), .B (n_242), .Q (out_0[30]));
  EN2X1 g2713(.A (n_297), .B (n_241), .Q (out_0[29]));
  EN2X1 g2714(.A (n_295), .B (n_240), .Q (out_0[28]));
  EN2X1 g2715(.A (n_293), .B (n_239), .Q (out_0[27]));
  EN2X1 g2716(.A (n_280), .B (n_228), .Q (out_0[21]));
  EO2X1 g2717(.A (n_289), .B (n_227), .Q (out_0[25]));
  EO2X1 g2718(.A (n_301), .B (n_310), .Q (out_0[31]));
  NO2I1X4 g2723(.B (n_303), .AN (n_187), .Q (n_304));
  AN21X1 g3(.A (n_166), .B (n_288), .C (n_190), .Q (n_303));
  INX1 g2724(.A (n_305), .Q (n_306));
  NO3X2 g2726(.A (n_273), .B (n_191), .C (n_189), .Q (n_307));
  NA3X2 g2727(.A (n_257), .B (n_174), .C (n_173), .Q (n_308));
  EO3X1 g2728(.A (in_1[0]), .B (in_2[0]), .C (in_0[0]), .Q (out_0[0]));
  EN3X1 g2729(.A (in_1[31]), .B (in_0[31]), .C (n_153), .Q (n_310));
  HAX2 g2730(.A (in_1[4]), .B (in_0[4]), .S (n_312), .CO (n_311));
  FAX1 g2732(.A (in_1[0]), .B (in_2[0]), .CI (in_0[0]), .S
       (UNCONNECTED), .CO (n_305));
endmodule

module rvsteel_core(clock, reset, halt, rw_address, read_data,
     read_request, read_response, write_data, write_strobe,
     write_request, write_response, irq_external,
     irq_external_response, irq_timer, irq_timer_response,
     irq_software, irq_software_response, irq_fast, irq_fast_response,
     real_time_clock);
  input clock, reset, halt, read_response, write_response,
       irq_external, irq_timer, irq_software;
  input [31:0] read_data;
  input [15:0] irq_fast;
  input [63:0] real_time_clock;
  output [31:0] rw_address, write_data;
  output read_request, write_request, irq_external_response,
       irq_timer_response, irq_software_response;
  output [3:0] write_strobe;
  output [15:0] irq_fast_response;
  wire clock, reset, halt, read_response, write_response, irq_external,
       irq_timer, irq_software;
  wire [31:0] read_data;
  wire [15:0] irq_fast;
  wire [63:0] real_time_clock;
  wire [31:0] rw_address, write_data;
  wire read_request, write_request, irq_external_response,
       irq_timer_response, irq_software_response;
  wire [3:0] write_strobe;
  wire [15:0] irq_fast_response;
  wire [31:0] alu_sra_result;
  wire [31:0] alu_2nd_operand;
  wire [3:0] current_state;
  wire [31:0] instruction;
  wire [31:0] prev_instruction;
  wire [63:0] csr_utime;
  wire [31:0] instruction_address;
  wire [31:0] prev_rw_address;
  wire [31:0] csr_data_out;
  wire [63:0] csr_minstret;
  wire [63:0] csr_mcycle;
  wire [31:0] prev_instruction_address;
  wire [31:0] csr_mcause;
  wire [31:0] csr_mtval;
  wire [31:0] csr_mscratch;
  wire [3:0] prev_write_strobe;
  wire [31:0] program_counter;
  wire [31:0] prev_write_data;
  wire [31:0] csr_mtvec;
  wire [4:0] csr_mcause_code;
  wire UNCONNECTED_HIER_Z, UNCONNECTED_HIER_Z0, UNCONNECTED_HIER_Z1,
       UNCONNECTED_HIER_Z2, UNCONNECTED_HIER_Z3, UNCONNECTED_HIER_Z4,
       UNCONNECTED_HIER_Z5, UNCONNECTED_HIER_Z6;
  wire UNCONNECTED_HIER_Z7, UNCONNECTED_HIER_Z8, UNCONNECTED_HIER_Z9,
       UNCONNECTED_HIER_Z10, UNCONNECTED_HIER_Z11,
       UNCONNECTED_HIER_Z12, UNCONNECTED_HIER_Z13, UNCONNECTED_HIER_Z14;
  wire UNCONNECTED_HIER_Z15, UNCONNECTED_HIER_Z16,
       UNCONNECTED_HIER_Z17, UNCONNECTED_HIER_Z18,
       UNCONNECTED_HIER_Z19, UNCONNECTED_HIER_Z20,
       UNCONNECTED_HIER_Z21, UNCONNECTED_HIER_Z22;
  wire UNCONNECTED_HIER_Z23, UNCONNECTED_HIER_Z24,
       UNCONNECTED_HIER_Z25, UNCONNECTED_HIER_Z26,
       UNCONNECTED_HIER_Z27, UNCONNECTED_HIER_Z28,
       UNCONNECTED_HIER_Z29, UNCONNECTED_HIER_Z30;
  wire UNCONNECTED_HIER_Z31, UNCONNECTED_HIER_Z32,
       UNCONNECTED_HIER_Z33, add_459_21_n_755, add_459_21_n_758,
       add_459_21_n_761, add_459_21_n_764, add_459_21_n_766;
  wire add_459_21_n_769, add_459_21_n_771, add_459_21_n_774,
       add_459_21_n_776, add_459_21_n_778, add_459_21_n_780,
       add_459_21_n_782, add_459_21_n_784;
  wire add_459_21_n_786, add_459_21_n_788, add_459_21_n_790,
       add_459_21_n_792, add_459_21_n_794, add_459_21_n_795,
       add_459_21_n_802, add_459_21_n_803;
  wire add_459_21_n_810, add_459_21_n_811, add_459_21_n_818,
       add_459_21_n_819, add_459_21_n_825, add_459_21_n_831,
       add_459_21_n_837, add_463_14_n_598;
  wire add_463_14_n_601, add_463_14_n_603, add_463_14_n_608,
       add_463_14_n_610, add_463_14_n_613, add_463_14_n_614,
       add_463_14_n_615, add_463_14_n_618;
  wire add_463_14_n_620, add_463_14_n_629, add_463_14_n_631,
       add_463_14_n_633, add_463_14_n_635, add_463_14_n_636,
       add_463_14_n_639, add_463_14_n_640;
  wire add_463_14_n_644, add_463_14_n_647, add_463_14_n_648,
       add_463_14_n_650, add_463_14_n_653, add_463_14_n_654,
       add_463_14_n_655, add_463_14_n_662;
  wire add_463_14_n_663, add_463_14_n_664, add_463_14_n_667,
       add_463_14_n_669, add_463_14_n_673, add_463_14_n_676,
       add_463_14_n_679, add_463_14_n_683;
  wire add_463_14_n_685, add_463_14_n_687, add_463_14_n_688,
       add_463_14_n_691, add_463_14_n_694, add_463_14_n_695,
       add_463_14_n_696, add_463_14_n_698;
  wire add_463_14_n_700, add_463_14_n_702, add_463_14_n_705,
       add_463_14_n_706, add_463_14_n_708, add_463_14_n_710,
       add_463_14_n_712, add_463_14_n_714;
  wire add_463_14_n_716, add_463_14_n_717, add_463_14_n_719,
       add_463_14_n_720, add_463_14_n_721, add_463_14_n_722,
       add_463_14_n_723, add_463_14_n_724;
  wire add_463_14_n_725, add_463_14_n_726, add_463_14_n_727,
       add_463_14_n_728, add_463_14_n_738, add_463_14_n_739,
       add_463_14_n_740, add_463_14_n_741;
  wire add_463_14_n_742, add_463_14_n_743, add_463_14_n_744,
       add_463_14_n_748, add_463_14_n_756, add_463_14_n_757,
       add_463_14_n_758, add_463_14_n_759;
  wire add_463_14_n_760, add_463_14_n_761, add_463_14_n_762,
       add_463_14_n_763, add_463_14_n_764, add_463_14_n_765,
       add_463_14_n_766, add_463_14_n_771;
  wire add_463_14_n_774, add_463_14_n_776, add_463_14_n_780,
       add_463_14_n_782, add_463_14_n_784, add_463_14_n_785,
       add_463_14_n_788, add_463_14_n_789;
  wire add_463_14_n_791, add_463_14_n_795, add_463_14_n_796,
       add_463_14_n_798, add_463_14_n_800, add_463_14_n_802,
       add_463_14_n_803, add_463_14_n_805;
  wire add_463_14_n_807, add_463_14_n_808, add_463_14_n_809,
       add_463_14_n_810, add_463_14_n_811, add_463_14_n_812,
       add_463_14_n_814, add_463_14_n_816;
  wire add_463_14_n_817, add_463_14_n_819, add_463_14_n_821,
       add_463_14_n_824, add_463_14_n_826, add_463_14_n_829,
       add_463_14_n_830, add_463_14_n_831;
  wire add_463_14_n_832, add_463_14_n_833, add_463_14_n_834,
       add_463_14_n_835, add_463_14_n_836, add_463_14_n_837,
       add_463_14_n_838, add_463_14_n_839;
  wire add_463_14_n_840, add_463_14_n_841, add_463_14_n_842,
       add_463_14_n_843, add_463_14_n_844, add_463_14_n_845,
       add_463_14_n_846, add_463_14_n_847;
  wire add_463_14_n_848, add_463_14_n_849, add_463_14_n_850,
       add_463_14_n_851, add_463_14_n_852, add_463_14_n_853,
       add_463_14_n_854, add_463_14_n_855;
  wire add_463_14_n_856, add_463_14_n_857, add_463_14_n_858,
       add_463_14_n_877, add_463_14_n_878, add_463_14_n_879,
       add_463_14_n_880, add_463_14_n_881;
  wire add_463_14_n_882, add_463_14_n_883, add_463_14_n_884,
       add_463_14_n_885, add_463_14_n_886, add_463_14_n_887,
       add_463_14_n_888, add_463_14_n_889;
  wire add_463_14_n_890, add_463_14_n_891, add_463_14_n_892,
       add_463_14_n_893, add_463_14_n_894, add_463_14_n_895,
       add_463_14_n_896, add_463_14_n_897;
  wire add_463_14_n_898, add_463_14_n_899, add_463_14_n_900,
       add_463_14_n_901, add_463_14_n_902, add_463_14_n_903,
       add_463_14_n_904, add_463_14_n_905;
  wire add_463_14_n_906, add_463_14_n_937, add_464_21_n_598,
       add_464_21_n_600, add_464_21_n_603, add_464_21_n_607,
       add_464_21_n_610, add_464_21_n_613;
  wire add_464_21_n_614, add_464_21_n_616, add_464_21_n_618,
       add_464_21_n_620, add_464_21_n_623, add_464_21_n_624,
       add_464_21_n_626, add_464_21_n_628;
  wire add_464_21_n_631, add_464_21_n_639, add_464_21_n_640,
       add_464_21_n_641, add_464_21_n_644, add_464_21_n_650,
       add_464_21_n_652, add_464_21_n_656;
  wire add_464_21_n_659, add_464_21_n_662, add_464_21_n_663,
       add_464_21_n_665, add_464_21_n_666, add_464_21_n_669,
       add_464_21_n_673, add_464_21_n_674;
  wire add_464_21_n_676, add_464_21_n_680, add_464_21_n_681,
       add_464_21_n_684, add_464_21_n_687, add_464_21_n_690,
       add_464_21_n_691, add_464_21_n_692;
  wire add_464_21_n_695, add_464_21_n_697, add_464_21_n_699,
       add_464_21_n_700, add_464_21_n_702, add_464_21_n_703,
       add_464_21_n_705, add_464_21_n_707;
  wire add_464_21_n_709, add_464_21_n_711, add_464_21_n_712,
       add_464_21_n_714, add_464_21_n_716, add_464_21_n_718,
       add_464_21_n_720, add_464_21_n_721;
  wire add_464_21_n_722, add_464_21_n_723, add_464_21_n_724,
       add_464_21_n_725, add_464_21_n_726, add_464_21_n_727,
       add_464_21_n_728, add_464_21_n_729;
  wire add_464_21_n_731, add_464_21_n_740, add_464_21_n_741,
       add_464_21_n_742, add_464_21_n_743, add_464_21_n_744,
       add_464_21_n_745, add_464_21_n_746;
  wire add_464_21_n_747, add_464_21_n_748, add_464_21_n_756,
       add_464_21_n_757, add_464_21_n_758, add_464_21_n_759,
       add_464_21_n_760, add_464_21_n_761;
  wire add_464_21_n_762, add_464_21_n_763, add_464_21_n_768,
       add_464_21_n_770, add_464_21_n_771, add_464_21_n_773,
       add_464_21_n_775, add_464_21_n_777;
  wire add_464_21_n_780, add_464_21_n_782, add_464_21_n_783,
       add_464_21_n_785, add_464_21_n_786, add_464_21_n_789,
       add_464_21_n_792, add_464_21_n_795;
  wire add_464_21_n_796, add_464_21_n_797, add_464_21_n_798,
       add_464_21_n_799, add_464_21_n_800, add_464_21_n_802,
       add_464_21_n_803, add_464_21_n_805;
  wire add_464_21_n_808, add_464_21_n_809, add_464_21_n_810,
       add_464_21_n_813, add_464_21_n_815, add_464_21_n_816,
       add_464_21_n_819, add_464_21_n_821;
  wire add_464_21_n_824, add_464_21_n_827, add_464_21_n_829,
       add_464_21_n_830, add_464_21_n_832, add_464_21_n_833,
       add_464_21_n_834, add_464_21_n_835;
  wire add_464_21_n_836, add_464_21_n_837, add_464_21_n_838,
       add_464_21_n_839, add_464_21_n_840, add_464_21_n_841,
       add_464_21_n_842, add_464_21_n_843;
  wire add_464_21_n_844, add_464_21_n_845, add_464_21_n_846,
       add_464_21_n_847, add_464_21_n_848, add_464_21_n_849,
       add_464_21_n_850, add_464_21_n_851;
  wire add_464_21_n_852, add_464_21_n_853, add_464_21_n_854,
       add_464_21_n_855, add_464_21_n_856, add_464_21_n_857,
       add_464_21_n_858, add_464_21_n_859;
  wire add_464_21_n_860, add_464_21_n_861, add_464_21_n_890,
       add_464_21_n_891, add_464_21_n_892, add_464_21_n_893,
       add_464_21_n_894, add_464_21_n_895;
  wire add_464_21_n_896, add_464_21_n_897, add_464_21_n_898,
       add_464_21_n_899, add_464_21_n_900, add_464_21_n_901,
       add_464_21_n_902, add_464_21_n_903;
  wire add_464_21_n_904, add_464_21_n_905, add_464_21_n_906,
       add_464_21_n_907, add_464_21_n_908, add_464_21_n_909,
       add_464_21_n_910, add_464_21_n_911;
  wire add_464_21_n_912, add_464_21_n_913, add_464_21_n_914,
       add_464_21_n_915, add_464_21_n_916, add_464_21_n_917,
       add_464_21_n_918, add_464_21_n_919;
  wire add_464_21_n_920, add_1545_30_n_700, add_1545_30_n_703,
       add_1545_30_n_706, add_1545_30_n_710, add_1545_30_n_712,
       add_1545_30_n_715, add_1545_30_n_717;
  wire add_1545_30_n_719, add_1545_30_n_721, add_1545_30_n_723,
       add_1545_30_n_725, add_1545_30_n_727, add_1545_30_n_729,
       add_1545_30_n_731, add_1545_30_n_732;
  wire add_1545_30_n_737, add_1545_30_n_738, add_1545_30_n_745,
       add_1545_30_n_746, add_1545_30_n_753, add_1545_30_n_754,
       add_1545_30_n_760, add_1545_30_n_766;
  wire add_1545_30_n_772, add_1545_30_n_775, add_1545_30_n_777,
       add_1545_30_n_779, add_1545_30_n_781, add_1545_30_n_783,
       alu_operation_code_39061, branch_type;
  wire csr_mcause_interrupt_flag, flush_37507,
       inc_ADD_UNS_OP5493_6_n_452, inc_ADD_UNS_OP5493_6_n_454,
       inc_ADD_UNS_OP5493_6_n_456, inc_ADD_UNS_OP5493_6_n_458,
       inc_ADD_UNS_OP5493_6_n_460, inc_ADD_UNS_OP5493_6_n_462;
  wire inc_ADD_UNS_OP5493_6_n_464, inc_ADD_UNS_OP5493_6_n_466,
       inc_ADD_UNS_OP5493_6_n_468, inc_ADD_UNS_OP5493_6_n_470,
       inc_ADD_UNS_OP5493_6_n_472, inc_ADD_UNS_OP5493_6_n_474,
       inc_ADD_UNS_OP5493_6_n_483, inc_ADD_UNS_OP5493_6_n_488;
  wire inc_ADD_UNS_OP5493_6_n_493, inc_ADD_UNS_OP5493_6_n_498,
       inc_ADD_UNS_OP5493_6_n_503, inc_ADD_UNS_OP5493_6_n_508,
       inc_ADD_UNS_OP5493_6_n_511, inc_ADD_UNS_OP5493_6_n_514,
       inc_ADD_UNS_OP5493_6_n_517, inc_ADD_UNS_OP5493_6_n_520;
  wire inc_ADD_UNS_OP5493_6_n_525, inc_ADD_UNS_OP5493_6_n_528,
       inc_ADD_UNS_OP5493_6_n_531, inc_ADD_UNS_OP5493_6_n_534,
       inc_ADD_UNS_OP5493_6_n_537, inc_ADD_UNS_OP5493_6_n_540,
       inc_ADD_UNS_OP5493_6_n_542, inc_ADD_UNS_OP5493_6_n_545;
  wire inc_ADD_UNS_OP5493_6_n_550, inc_ADD_UNS_OP5493_6_n_553,
       inc_ADD_UNS_OP5493_6_n_558, inc_ADD_UNS_OP5493_6_n_563,
       inc_ADD_UNS_OP5493_6_n_568, inc_ADD_UNS_OP5493_6_n_571,
       inc_ADD_UNS_OP5493_6_n_576, inc_ADD_UNS_OP5493_6_n_581;
  wire inc_ADD_UNS_OP5493_6_n_586, inc_ADD_UNS_OP5493_6_n_591,
       inc_ADD_UNS_OP5493_6_n_594, inc_ADD_UNS_OP5493_6_n_599,
       inc_ADD_UNS_OP5493_6_n_602, inc_ADD_UNS_OP5493_6_n_607,
       inc_ADD_UNS_OP5493_6_n_610, inc_ADD_UNS_OP5493_6_n_613;
  wire inc_ADD_UNS_OP5493_6_n_616, inc_ADD_UNS_OP5493_6_n_619,
       inc_ADD_UNS_OP5493_6_n_622, inc_ADD_UNS_OP5493_6_n_625,
       inc_ADD_UNS_OP5493_6_n_630, inc_ADD_UNS_OP5493_6_n_635,
       inc_ADD_UNS_OP5493_6_n_650, inc_ADD_UNS_OP5493_6_n_655;
  wire inc_ADD_UNS_OP5493_6_n_660, inc_ADD_UNS_OP5493_6_n_665,
       inc_ADD_UNS_OP5493_6_n_668, inc_ADD_UNS_OP5493_6_n_671,
       inc_ADD_UNS_OP5493_6_n_674, inc_ADD_UNS_OP5493_6_n_677,
       inc_ADD_UNS_OP5493_6_n_737, inc_ADD_UNS_OP5493_6_n_738;
  wire inc_ADD_UNS_OP5493_6_n_741, inc_ADD_UNS_OP5494_3_n_452,
       inc_ADD_UNS_OP5494_3_n_455, inc_ADD_UNS_OP5494_3_n_458,
       inc_ADD_UNS_OP5494_3_n_460, inc_ADD_UNS_OP5494_3_n_462,
       inc_ADD_UNS_OP5494_3_n_464, inc_ADD_UNS_OP5494_3_n_466;
  wire inc_ADD_UNS_OP5494_3_n_468, inc_ADD_UNS_OP5494_3_n_470,
       inc_ADD_UNS_OP5494_3_n_472, inc_ADD_UNS_OP5494_3_n_474,
       inc_ADD_UNS_OP5494_3_n_476, inc_ADD_UNS_OP5494_3_n_478,
       inc_ADD_UNS_OP5494_3_n_483, inc_ADD_UNS_OP5494_3_n_488;
  wire inc_ADD_UNS_OP5494_3_n_493, inc_ADD_UNS_OP5494_3_n_498,
       inc_ADD_UNS_OP5494_3_n_503, inc_ADD_UNS_OP5494_3_n_508,
       inc_ADD_UNS_OP5494_3_n_513, inc_ADD_UNS_OP5494_3_n_518,
       inc_ADD_UNS_OP5494_3_n_521, inc_ADD_UNS_OP5494_3_n_524;
  wire inc_ADD_UNS_OP5494_3_n_527, inc_ADD_UNS_OP5494_3_n_530,
       inc_ADD_UNS_OP5494_3_n_533, inc_ADD_UNS_OP5494_3_n_536,
       inc_ADD_UNS_OP5494_3_n_539, inc_ADD_UNS_OP5494_3_n_542,
       inc_ADD_UNS_OP5494_3_n_545, inc_ADD_UNS_OP5494_3_n_548;
  wire inc_ADD_UNS_OP5494_3_n_551, inc_ADD_UNS_OP5494_3_n_554,
       inc_ADD_UNS_OP5494_3_n_557, inc_ADD_UNS_OP5494_3_n_562,
       inc_ADD_UNS_OP5494_3_n_567, inc_ADD_UNS_OP5494_3_n_572,
       inc_ADD_UNS_OP5494_3_n_577, inc_ADD_UNS_OP5494_3_n_582;
  wire inc_ADD_UNS_OP5494_3_n_585, inc_ADD_UNS_OP5494_3_n_588,
       inc_ADD_UNS_OP5494_3_n_591, inc_ADD_UNS_OP5494_3_n_594,
       inc_ADD_UNS_OP5494_3_n_599, inc_ADD_UNS_OP5494_3_n_604,
       inc_ADD_UNS_OP5494_3_n_607, inc_ADD_UNS_OP5494_3_n_610;
  wire inc_ADD_UNS_OP5494_3_n_613, inc_ADD_UNS_OP5494_3_n_616,
       inc_ADD_UNS_OP5494_3_n_631, inc_ADD_UNS_OP5494_3_n_636,
       inc_ADD_UNS_OP5494_3_n_641, inc_ADD_UNS_OP5494_3_n_646,
       inc_ADD_UNS_OP5494_3_n_651, inc_ADD_UNS_OP5494_3_n_661;
  wire inc_ADD_UNS_OP5494_3_n_664, inc_ADD_UNS_OP5494_3_n_667,
       inc_ADD_UNS_OP5494_3_n_670, inc_ADD_UNS_OP5494_3_n_673,
       inc_ADD_UNS_OP5494_3_n_676, inc_ADD_UNS_OP5494_3_n_736,
       inc_ADD_UNS_OP5494_3_n_737, inc_ADD_UNS_OP5494_3_n_740;
  wire inc_ADD_UNS_OP_5_n_2648, inc_ADD_UNS_OP_5_n_2652,
       inc_ADD_UNS_OP_5_n_2656, inc_ADD_UNS_OP_5_n_2661,
       inc_ADD_UNS_OP_5_n_2665, inc_ADD_UNS_OP_5_n_2667,
       inc_ADD_UNS_OP_5_n_2672, inc_ADD_UNS_OP_5_n_2678;
  wire inc_ADD_UNS_OP_5_n_2683, inc_ADD_UNS_OP_5_n_2688,
       inc_ADD_UNS_OP_5_n_2693, inc_ADD_UNS_OP_5_n_2699,
       inc_ADD_UNS_OP_5_n_2704, inc_ADD_UNS_OP_5_n_2708,
       inc_ADD_UNS_OP_5_n_2710, inc_ADD_UNS_OP_5_n_2718;
  wire inc_ADD_UNS_OP_5_n_2720, inc_ADD_UNS_OP_5_n_2724,
       inc_ADD_UNS_OP_5_n_2727, inc_ADD_UNS_OP_5_n_2730,
       inc_ADD_UNS_OP_5_n_2738, inc_ADD_UNS_OP_5_n_2740,
       inc_ADD_UNS_OP_5_n_2744, inc_ADD_UNS_OP_5_n_2747;
  wire inc_ADD_UNS_OP_5_n_2752, inc_ADD_UNS_OP_5_n_2756,
       inc_ADD_UNS_OP_5_n_2758, inc_ADD_UNS_OP_5_n_2762,
       inc_ADD_UNS_OP_5_n_2765, inc_ADD_UNS_OP_5_n_2770,
       inc_ADD_UNS_OP_5_n_2774, inc_ADD_UNS_OP_5_n_2776;
  wire inc_ADD_UNS_OP_5_n_2780, inc_ADD_UNS_OP_5_n_2783,
       inc_ADD_UNS_OP_5_n_2788, inc_ADD_UNS_OP_5_n_2791,
       inc_ADD_UNS_OP_5_n_2794, inc_ADD_UNS_OP_5_n_2797,
       inc_ADD_UNS_OP_5_n_2800, inc_ADD_UNS_OP_5_n_2805;
  wire inc_ADD_UNS_OP_5_n_2808, inc_ADD_UNS_OP_5_n_2811,
       inc_ADD_UNS_OP_5_n_2814, inc_ADD_UNS_OP_5_n_2817,
       inc_ADD_UNS_OP_5_n_2820, inc_ADD_UNS_OP_5_n_2823,
       inc_ADD_UNS_OP_5_n_2825, inc_ADD_UNS_OP_5_n_2828;
  wire inc_ADD_UNS_OP_5_n_2831, inc_ADD_UNS_OP_5_n_2834,
       inc_ADD_UNS_OP_5_n_2837, inc_ADD_UNS_OP_5_n_2840,
       inc_ADD_UNS_OP_5_n_2842, inc_ADD_UNS_OP_5_n_2844,
       inc_ADD_UNS_OP_5_n_2847, inc_ADD_UNS_OP_5_n_2850;
  wire inc_ADD_UNS_OP_5_n_2855, inc_ADD_UNS_OP_5_n_2860,
       inc_ADD_UNS_OP_5_n_2868, inc_ADD_UNS_OP_5_n_2871,
       inc_ADD_UNS_OP_5_n_2876, inc_ADD_UNS_OP_5_n_2881,
       inc_ADD_UNS_OP_5_n_2886, inc_ADD_UNS_OP_5_n_2889;
  wire inc_ADD_UNS_OP_5_n_2891, inc_ADD_UNS_OP_5_n_2894,
       inc_ADD_UNS_OP_5_n_2924, inc_ADD_UNS_OP_5_n_2929,
       inc_ADD_UNS_OP_5_n_2931, inc_ADD_UNS_OP_5_n_2948,
       inc_ADD_UNS_OP_5_n_2966, inc_ADD_UNS_OP_5_n_2968;
  wire inc_ADD_UNS_OP_5_n_2970, inc_ADD_UNS_OP_5_n_2973,
       inc_ADD_UNS_OP_5_n_2974, inc_ADD_UNS_OP_5_n_2987,
       inc_add_1343_59_4_n_703, inc_add_1343_59_4_n_708,
       inc_add_1343_59_4_n_713, inc_add_1343_59_4_n_718;
  wire inc_add_1343_59_4_n_724, inc_add_1343_59_4_n_727,
       inc_add_1343_59_4_n_735, inc_add_1343_59_4_n_740,
       inc_add_1343_59_4_n_745, inc_add_1343_59_4_n_751,
       inc_add_1343_59_4_n_753, inc_add_1343_59_4_n_758;
  wire inc_add_1343_59_4_n_761, inc_add_1343_59_4_n_763,
       inc_add_1343_59_4_n_771, inc_add_1343_59_4_n_773,
       inc_add_1343_59_4_n_777, inc_add_1343_59_4_n_780,
       inc_add_1343_59_4_n_783, inc_add_1343_59_4_n_791;
  wire inc_add_1343_59_4_n_793, inc_add_1343_59_4_n_797,
       inc_add_1343_59_4_n_800, inc_add_1343_59_4_n_805,
       inc_add_1343_59_4_n_809, inc_add_1343_59_4_n_811,
       inc_add_1343_59_4_n_815, inc_add_1343_59_4_n_819;
  wire inc_add_1343_59_4_n_824, inc_add_1343_59_4_n_830,
       inc_add_1343_59_4_n_832, inc_add_1343_59_4_n_834,
       inc_add_1343_59_4_n_835, inc_add_1343_59_4_n_841,
       inc_add_1343_59_4_n_844, inc_add_1343_59_4_n_847;
  wire inc_add_1343_59_4_n_850, inc_add_1343_59_4_n_855,
       inc_add_1343_59_4_n_858, inc_add_1343_59_4_n_861,
       inc_add_1343_59_4_n_864, inc_add_1343_59_4_n_867,
       inc_add_1343_59_4_n_870, inc_add_1343_59_4_n_873;
  wire inc_add_1343_59_4_n_876, inc_add_1343_59_4_n_879,
       inc_add_1343_59_4_n_882, inc_add_1343_59_4_n_885,
       inc_add_1343_59_4_n_888, inc_add_1343_59_4_n_890,
       inc_add_1343_59_4_n_892, inc_add_1343_59_4_n_894;
  wire inc_add_1343_59_4_n_896, inc_add_1343_59_4_n_898,
       inc_add_1343_59_4_n_900, inc_add_1343_59_4_n_905,
       inc_add_1343_59_4_n_911, inc_add_1343_59_4_n_914,
       inc_add_1343_59_4_n_918, inc_add_1343_59_4_n_923;
  wire inc_add_1343_59_4_n_925, inc_add_1343_59_4_n_929,
       inc_add_1343_59_4_n_930, inc_add_1343_59_4_n_968,
       inc_add_1343_59_4_n_972, inc_add_1343_59_4_n_992,
       inc_add_1343_59_4_n_1007, inc_add_1343_59_4_n_1010;
  wire inc_add_1345_58_1_n_448, inc_add_1345_58_1_n_451,
       inc_add_1345_58_1_n_454, inc_add_1345_58_1_n_456,
       inc_add_1345_58_1_n_458, inc_add_1345_58_1_n_460,
       inc_add_1345_58_1_n_462, inc_add_1345_58_1_n_464;
  wire inc_add_1345_58_1_n_466, inc_add_1345_58_1_n_471,
       inc_add_1345_58_1_n_476, inc_add_1345_58_1_n_481,
       inc_add_1345_58_1_n_486, inc_add_1345_58_1_n_494,
       inc_add_1345_58_1_n_497, inc_add_1345_58_1_n_499;
  wire inc_add_1345_58_1_n_504, inc_add_1345_58_1_n_509,
       inc_add_1345_58_1_n_514, inc_add_1345_58_1_n_517,
       inc_add_1345_58_1_n_520, inc_add_1345_58_1_n_525,
       inc_add_1345_58_1_n_528, inc_add_1345_58_1_n_531;
  wire inc_add_1345_58_1_n_534, inc_add_1345_58_1_n_537,
       inc_add_1345_58_1_n_539, inc_add_1345_58_1_n_544,
       inc_add_1345_58_1_n_547, inc_add_1345_58_1_n_550,
       inc_add_1345_58_1_n_553, inc_add_1345_58_1_n_556;
  wire inc_add_1345_58_1_n_559, inc_add_1345_58_1_n_562,
       inc_add_1345_58_1_n_565, inc_add_1345_58_1_n_568,
       inc_add_1345_58_1_n_573, inc_add_1345_58_1_n_576,
       inc_add_1345_58_1_n_579, inc_add_1345_58_1_n_582;
  wire inc_add_1345_58_1_n_585, inc_add_1345_58_1_n_590,
       inc_add_1345_58_1_n_595, inc_add_1345_58_1_n_600,
       inc_add_1345_58_1_n_605, inc_add_1345_58_1_n_608,
       inc_add_1345_58_1_n_611, inc_add_1345_58_1_n_614;
  wire inc_add_1345_58_1_n_617, inc_add_1345_58_1_n_627,
       inc_add_1345_58_1_n_630, inc_add_1345_58_1_n_633,
       inc_add_1345_58_1_n_638, inc_add_1345_58_1_n_643,
       inc_add_1345_58_1_n_648, inc_add_1345_58_1_n_653;
  wire inc_add_1345_58_1_n_658, inc_add_1345_58_1_n_663,
       inc_add_1345_58_1_n_668, inc_add_1345_58_1_n_673,
       inc_add_1345_58_1_n_728, inc_add_1345_58_1_n_732,
       inc_add_1347_34_2_n_448, inc_add_1347_34_2_n_451;
  wire inc_add_1347_34_2_n_454, inc_add_1347_34_2_n_456,
       inc_add_1347_34_2_n_458, inc_add_1347_34_2_n_460,
       inc_add_1347_34_2_n_462, inc_add_1347_34_2_n_464,
       inc_add_1347_34_2_n_466, inc_add_1347_34_2_n_468;
  wire inc_add_1347_34_2_n_470, inc_add_1347_34_2_n_472,
       inc_add_1347_34_2_n_474, inc_add_1347_34_2_n_479,
       inc_add_1347_34_2_n_484, inc_add_1347_34_2_n_489,
       inc_add_1347_34_2_n_494, inc_add_1347_34_2_n_499;
  wire inc_add_1347_34_2_n_504, inc_add_1347_34_2_n_509,
       inc_add_1347_34_2_n_514, inc_add_1347_34_2_n_517,
       inc_add_1347_34_2_n_520, inc_add_1347_34_2_n_523,
       inc_add_1347_34_2_n_526, inc_add_1347_34_2_n_529;
  wire inc_add_1347_34_2_n_532, inc_add_1347_34_2_n_535,
       inc_add_1347_34_2_n_538, inc_add_1347_34_2_n_541,
       inc_add_1347_34_2_n_546, inc_add_1347_34_2_n_549,
       inc_add_1347_34_2_n_552, inc_add_1347_34_2_n_555;
  wire inc_add_1347_34_2_n_558, inc_add_1347_34_2_n_563,
       inc_add_1347_34_2_n_568, inc_add_1347_34_2_n_571,
       inc_add_1347_34_2_n_574, inc_add_1347_34_2_n_577,
       inc_add_1347_34_2_n_580, inc_add_1347_34_2_n_585;
  wire inc_add_1347_34_2_n_590, inc_add_1347_34_2_n_595,
       inc_add_1347_34_2_n_598, inc_add_1347_34_2_n_601,
       inc_add_1347_34_2_n_604, inc_add_1347_34_2_n_607,
       inc_add_1347_34_2_n_612, inc_add_1347_34_2_n_617;
  wire inc_add_1347_34_2_n_620, inc_add_1347_34_2_n_623,
       inc_add_1347_34_2_n_626, inc_add_1347_34_2_n_629,
       inc_add_1347_34_2_n_634, inc_add_1347_34_2_n_639,
       inc_add_1347_34_2_n_644, inc_add_1347_34_2_n_649;
  wire inc_add_1347_34_2_n_654, inc_add_1347_34_2_n_659,
       inc_add_1347_34_2_n_664, inc_add_1347_34_2_n_669,
       \instruction[5]_40139 , \instruction[7]_39562 ,
       \instruction[8]_40015 , \instruction[9]_39983 ;
  wire \instruction[10]_39951 , \instruction[11]_40800 ,
       \instruction[14]_40077 , jal_type, jalr_type, load_request_BAR,
       mret, n_0;
  wire n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_9;
  wire n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17;
  wire n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25;
  wire n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33;
  wire n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41;
  wire n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666;
  wire n_667, n_668, n_669, n_670, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_678, n_679, n_681, n_682, n_683, n_684;
  wire n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700;
  wire n_701, n_702, n_703, n_704, n_705, n_709, n_710, n_711;
  wire n_712, n_713, n_714, n_715, n_716, n_717, n_718, n_719;
  wire n_720, n_721, n_722, n_723, n_724, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760;
  wire n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784;
  wire n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792;
  wire n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800;
  wire n_801, n_802, n_803, n_804, n_805, n_806, n_807, n_808;
  wire n_809, n_811, n_812, n_814, n_815, n_816, n_817, n_818;
  wire n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826;
  wire n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834;
  wire n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842;
  wire n_843, n_844, n_845, n_846, n_848, n_849, n_850, n_851;
  wire n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859;
  wire n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867;
  wire n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875;
  wire n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883;
  wire n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891;
  wire n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899;
  wire n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907;
  wire n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956;
  wire n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964;
  wire n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972;
  wire n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980;
  wire n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988;
  wire n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996;
  wire n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004;
  wire n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012;
  wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028;
  wire n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036;
  wire n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044;
  wire n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052;
  wire n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060;
  wire n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068;
  wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084;
  wire n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092;
  wire n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100;
  wire n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108;
  wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116;
  wire n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124;
  wire n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132;
  wire n_1133, n_1134, n_1141, n_1142, n_1143, n_1144, n_1147, n_1148;
  wire n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156;
  wire n_1157, n_1159, n_1160, n_1161, n_1162, n_1163, n_1165, n_1166;
  wire n_1167, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175;
  wire n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183;
  wire n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191;
  wire n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207;
  wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
  wire n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223;
  wire n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231;
  wire n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239;
  wire n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247;
  wire n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255;
  wire n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263;
  wire n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271;
  wire n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279;
  wire n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287;
  wire n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295;
  wire n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303;
  wire n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311;
  wire n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319;
  wire n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327;
  wire n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335;
  wire n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343;
  wire n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351;
  wire n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359;
  wire n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367;
  wire n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375;
  wire n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383;
  wire n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391;
  wire n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399;
  wire n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407;
  wire n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415;
  wire n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423;
  wire n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431;
  wire n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439;
  wire n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447;
  wire n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455;
  wire n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463;
  wire n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471;
  wire n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487;
  wire n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495;
  wire n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503;
  wire n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511;
  wire n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519;
  wire n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527;
  wire n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535;
  wire n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543;
  wire n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551;
  wire n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567;
  wire n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575;
  wire n_1576, n_1577, n_1578, n_1580, n_1581, n_1582, n_1583, n_1584;
  wire n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592;
  wire n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601;
  wire n_1604, n_1605, n_1606, n_1608, n_1609, n_1611, n_1612, n_1613;
  wire n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621;
  wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629;
  wire n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637;
  wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645;
  wire n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653;
  wire n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1689, n_1690, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
  wire n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720;
  wire n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728;
  wire n_1729, n_1730, n_1731, n_1733, n_1734, n_1735, n_1736, n_1737;
  wire n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745;
  wire n_1746, n_1748, n_1750, n_1752, n_1753, n_1754, n_1755, n_1756;
  wire n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764;
  wire n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772;
  wire n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780;
  wire n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788;
  wire n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796;
  wire n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804;
  wire n_1805, n_1806, n_1807, n_1808, n_1809, n_1811, n_1812, n_1813;
  wire n_1814, n_1816, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1832, n_1833;
  wire n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841;
  wire n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849;
  wire n_1850, n_1851, n_1853, n_1854, n_1855, n_1856, n_1858, n_1859;
  wire n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867;
  wire n_1868, n_1869, n_1870, n_1872, n_1873, n_1874, n_1875, n_1876;
  wire n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886;
  wire n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894;
  wire n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902;
  wire n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910;
  wire n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918;
  wire n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926;
  wire n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934;
  wire n_1935, n_1936, n_1937, n_1938, n_1941, n_1942, n_1943, n_1944;
  wire n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960;
  wire n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976;
  wire n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984;
  wire n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992;
  wire n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000;
  wire n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008;
  wire n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016;
  wire n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024;
  wire n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032;
  wire n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040;
  wire n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048;
  wire n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056;
  wire n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064;
  wire n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072;
  wire n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080;
  wire n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088;
  wire n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096;
  wire n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104;
  wire n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112;
  wire n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120;
  wire n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128;
  wire n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136;
  wire n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144;
  wire n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152;
  wire n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160;
  wire n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168;
  wire n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176;
  wire n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184;
  wire n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192;
  wire n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200;
  wire n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208;
  wire n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216;
  wire n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224;
  wire n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232;
  wire n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240;
  wire n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248;
  wire n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256;
  wire n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264;
  wire n_2267, n_2268, n_2269, n_2270, n_2273, n_2274, n_2275, n_2276;
  wire n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284;
  wire n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292;
  wire n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300;
  wire n_2301, n_2302, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309;
  wire n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317;
  wire n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325;
  wire n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333;
  wire n_2334, n_2335, n_2336, n_2337, n_2338, n_2340, n_2341, n_2343;
  wire n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2353;
  wire n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2363;
  wire n_2364, n_2365, n_2366, n_2368, n_2369, n_2370, n_2371, n_2373;
  wire n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381;
  wire n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2390;
  wire n_2391, n_2393, n_2394, n_2395, n_2396, n_2398, n_2400, n_2401;
  wire n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409;
  wire n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2417, n_2418;
  wire n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426;
  wire n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434;
  wire n_2435, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452;
  wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460;
  wire n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468;
  wire n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476;
  wire n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484;
  wire n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492;
  wire n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500;
  wire n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508;
  wire n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516;
  wire n_2517, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525;
  wire n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533;
  wire n_2534, n_2535, n_2536, n_2537, n_2540, n_2541, n_2543, n_2544;
  wire n_2545, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553;
  wire n_2554, n_2555, n_2556, n_2557, n_2558, n_2560, n_2561, n_2563;
  wire n_2564, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2574;
  wire n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582;
  wire n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590;
  wire n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598;
  wire n_2599, n_2600, n_2601, n_2602, n_2603, n_2605, n_2606, n_2607;
  wire n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615;
  wire n_2616, n_2617, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624;
  wire n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632;
  wire n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640;
  wire n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648;
  wire n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656;
  wire n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664;
  wire n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672;
  wire n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680;
  wire n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688;
  wire n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696;
  wire n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704;
  wire n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712;
  wire n_2713, n_2714, n_2715, n_2716, n_2717, n_2719, n_2720, n_2721;
  wire n_2722, n_2723, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730;
  wire n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738;
  wire n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746;
  wire n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754;
  wire n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762;
  wire n_2763, n_2764, n_2765, n_2767, n_2768, n_2769, n_2770, n_2771;
  wire n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779;
  wire n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2788;
  wire n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796;
  wire n_2797, n_2798, n_2799, n_2800, n_2802, n_2803, n_2804, n_2805;
  wire n_2806, n_2807, n_2808, n_2811, n_2812, n_2813, n_2814, n_2815;
  wire n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2823, n_2824;
  wire n_2825, n_2826, n_2828, n_2829, n_2830, n_2833, n_2834, n_2835;
  wire n_2836, n_2838, n_2840, n_2842, n_2843, n_2844, n_2845, n_2846;
  wire n_2847, n_2848, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855;
  wire n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2863, n_2864;
  wire n_2865, n_2866, n_2867, n_2868, n_2869, n_2871, n_2872, n_2873;
  wire n_2874, n_2875, n_2878, n_2879, n_2881, n_2882, n_2883, n_2884;
  wire n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892;
  wire n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900;
  wire n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908;
  wire n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2918;
  wire n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926;
  wire n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934;
  wire n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942;
  wire n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950;
  wire n_2951, n_2952, n_2953, n_2955, n_2956, n_2959, n_2961, n_2962;
  wire n_2963, n_2965, n_2967, n_2969, n_2970, n_2971, n_2972, n_2973;
  wire n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981;
  wire n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989;
  wire n_2990, n_2992, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999;
  wire n_3000, n_3001, n_3002, n_3003, n_3005, n_3006, n_3007, n_3008;
  wire n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016;
  wire n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024;
  wire n_3025, n_3026, n_3027, n_3028, n_3030, n_3032, n_3033, n_3034;
  wire n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042;
  wire n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050;
  wire n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058;
  wire n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066;
  wire n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074;
  wire n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082;
  wire n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090;
  wire n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098;
  wire n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106;
  wire n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114;
  wire n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122;
  wire n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130;
  wire n_3131, n_3132, n_3133, n_3134, n_3135, n_3138, n_3139, n_3140;
  wire n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148;
  wire n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156;
  wire n_3157, n_3158, n_3160, n_3161, n_3162, n_3164, n_3166, n_3167;
  wire n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175;
  wire n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183;
  wire n_3184, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192;
  wire n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200;
  wire n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208;
  wire n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216;
  wire n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224;
  wire n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232;
  wire n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240;
  wire n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248;
  wire n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256;
  wire n_3257, n_3258, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265;
  wire n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273;
  wire n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281;
  wire n_3282, n_3283, n_3285, n_3287, n_3288, n_3290, n_3291, n_3292;
  wire n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300;
  wire n_3301, n_3302, n_3303, n_3304, n_3305, n_3309, n_3310, n_3311;
  wire n_3315, n_3316, n_3317, n_3318, n_3321, n_3322, n_3323, n_3324;
  wire n_3325, n_3326, n_3328, n_3329, n_3331, n_3332, n_3333, n_3334;
  wire n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342;
  wire n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350;
  wire n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358;
  wire n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366;
  wire n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374;
  wire n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382;
  wire n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390;
  wire n_3391, n_3392, n_3393, n_3394, n_3396, n_3397, n_3398, n_3399;
  wire n_3400, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408;
  wire n_3409, n_3410, n_3411, n_3414, n_3416, n_3420, n_3421, n_3422;
  wire n_3426, n_3428, n_3429, n_3430, n_3431, n_3433, n_3434, n_3435;
  wire n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, n_3443;
  wire n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451;
  wire n_3452, n_3453, n_3454, n_3455, n_3456, n_3458, n_3459, n_3460;
  wire n_3461, n_3462, n_3464, n_3465, n_3466, n_3467, n_3468, n_3471;
  wire n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479;
  wire n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487;
  wire n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495;
  wire n_3496, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504;
  wire n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512;
  wire n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520;
  wire n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528;
  wire n_3529, n_3530, n_3531, n_3534, n_3535, n_3536, n_3537, n_3538;
  wire n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546;
  wire n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554;
  wire n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564;
  wire n_3565, n_3566, n_3569, n_3570, n_3574, n_3575, n_3579, n_3580;
  wire n_3583, n_3586, n_3587, n_3588, n_3589, n_3592, n_3595, n_3599;
  wire n_3600, n_3603, n_3604, n_3607, n_3608, n_3609, n_3610, n_3611;
  wire n_3612, n_3613, n_3614, n_3617, n_3618, n_3619, n_3620, n_3621;
  wire n_3622, n_3625, n_3626, n_3633, n_3634, n_3649, n_3650, n_3653;
  wire n_3654, n_3657, n_3658, n_3663, n_3664, n_3665, n_3666, n_3667;
  wire n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675;
  wire n_3676, n_3677, n_3678, n_3681, n_3682, n_3683, n_3686, n_3687;
  wire n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, n_3695;
  wire n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703;
  wire n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711;
  wire n_3712, n_3713, n_3714, n_3715, n_3716, n_3719, n_3721, n_3724;
  wire n_3727, n_3728, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738;
  wire n_3739, n_3743, n_3744, n_3745, n_3747, n_3749, n_3750, n_3751;
  wire n_3752, n_3753, n_3754, n_3755, n_3758, n_3761, n_3762, n_3763;
  wire n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771;
  wire n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779;
  wire n_3780, n_3781, n_3782, n_3783, n_3784, n_3786, n_3787, n_3788;
  wire n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796;
  wire n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, n_3806, n_3807;
  wire n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815;
  wire n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823;
  wire n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831;
  wire n_3832, n_3834, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841;
  wire n_3843, n_3844, n_3845, n_3847, n_3850, n_3851, n_3852, n_3853;
  wire n_3854, n_3855, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863;
  wire n_3866, n_3868, n_3869, n_3871, n_3872, n_3874, n_3875, n_3877;
  wire n_3878, n_3879, n_3881, n_3882, n_3883, n_3884, n_3885, n_3886;
  wire n_3888, n_3890, n_3891, n_3893, n_3895, n_3897, n_3899, n_3900;
  wire n_3901, n_3902, n_3903, n_3904, n_3905, n_3907, n_3908, n_3909;
  wire n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3917, n_3919;
  wire n_3920, n_3923, n_3929, n_3930, n_3932, n_3935, n_3937, n_3938;
  wire n_3939, n_3942, n_3943, n_3944, n_3945, n_3946, n_3948, n_3949;
  wire n_3950, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958;
  wire n_3960, n_3962, n_3963, n_3965, n_3966, n_3967, n_3968, n_3969;
  wire n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978;
  wire n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986;
  wire n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994;
  wire n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001, n_4002;
  wire n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009, n_4010;
  wire n_4011, n_4012, n_4013, n_4014, n_4015, n_4017, n_4018, n_4019;
  wire n_4020, n_4021, n_4022, n_4023, n_4025, n_4026, n_4028, n_4030;
  wire n_4032, n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040;
  wire n_4041, n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048;
  wire n_4049, n_4050, n_4051, n_4052, n_4053, n_4055, n_4056, n_4057;
  wire n_4058, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066;
  wire n_4067, n_4069, n_4070, n_4071, n_4072, n_4073, n_4074, n_4075;
  wire n_4076, n_4078, n_4079, n_4080, n_4082, n_4083, n_4084, n_4085;
  wire n_4086, n_4087, n_4088, n_4090, n_4091, n_4092, n_4094, n_4098;
  wire n_4099, n_4101, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109;
  wire n_4110, n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117;
  wire n_4118, n_4119, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126;
  wire n_4127, n_4129, n_4130, n_4131, n_4132, n_4133, n_4135, n_4137;
  wire n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145;
  wire n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153;
  wire n_4154, n_4155, n_4156, n_4157, n_4159, n_4160, n_4161, n_4164;
  wire n_4165, n_4166, n_4167, n_4168, n_4169, n_4171, n_4172, n_4174;
  wire n_4175, n_4176, n_4177, n_4178, n_4179, n_4181, n_4183, n_4184;
  wire n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192;
  wire n_4194, n_4195, n_4196, n_4198, n_4199, n_4200, n_4202, n_4203;
  wire n_4204, n_4206, n_4207, n_4208, n_4209, n_4213, n_4215, n_4217;
  wire n_4218, n_4223, n_4227, n_4234, n_4235, n_4236, n_4239, n_4240;
  wire n_4241, n_4242, n_4243, n_4244, n_4245, n_4248, n_4249, n_4250;
  wire n_4251, n_4253, n_4258, n_4259, n_4260, n_4264, n_4265, n_4266;
  wire n_4267, n_4268, n_4275, n_4279, n_4280, n_4283, n_4284, n_4300;
  wire n_4301, n_4302, n_4303, n_4304, n_4307, n_4310, n_4311, n_4312;
  wire n_4313, n_4314, n_4315, n_4317, n_4320, n_4321, n_4322, n_4323;
  wire n_4324, n_4326, n_4328, n_4329, n_4330, n_4331, n_4333, n_4338;
  wire n_4343, n_4344, n_4352, n_4355, n_4356, n_4358, n_4360, n_4361;
  wire n_4362, n_4366, n_4367, n_4371, n_4372, n_4376, n_4377, n_4378;
  wire n_4379, n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386;
  wire n_4387, n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4396;
  wire n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403, n_4404;
  wire n_4405, n_4406, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415;
  wire n_4416, n_4417, n_4418, n_4419, n_4420, n_4422, n_4425, n_4426;
  wire n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4435, n_4436;
  wire n_4437, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445;
  wire n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4454, n_4455;
  wire n_4456, n_4457, n_4460, n_4461, n_4463, n_4464, n_4465, n_4466;
  wire n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481;
  wire n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4532, n_4533;
  wire n_4534, n_4535, n_4536, n_4538, n_4549, n_4550, n_4551, n_4552;
  wire n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560;
  wire n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568;
  wire n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576;
  wire n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584;
  wire n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592;
  wire n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600;
  wire n_4601, n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608;
  wire n_4609, n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616;
  wire n_4617, n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624;
  wire n_4625, n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632;
  wire n_4633, n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640;
  wire n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648;
  wire n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656;
  wire n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664;
  wire n_4665, n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672;
  wire n_4673, n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680;
  wire n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688;
  wire n_4689, n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696;
  wire n_4697, n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704;
  wire n_4705, n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712;
  wire n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720;
  wire n_4721, n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4728;
  wire n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735, n_4736;
  wire n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744;
  wire n_4745, n_4746, n_4747, n_4748, n_4749, n_4750, n_4751, n_4752;
  wire n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759, n_4760;
  wire n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767, n_4768;
  wire n_4769, n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776;
  wire n_4777, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784;
  wire n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4792;
  wire n_4793, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799, n_4800;
  wire n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808;
  wire n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816;
  wire n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824;
  wire n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832;
  wire n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840;
  wire n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4848;
  wire n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856;
  wire n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863, n_4864;
  wire n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872;
  wire n_4873, n_4874, n_4875, n_4876, n_4877, n_4878, n_4879, n_4880;
  wire n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888;
  wire n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896;
  wire n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4903, n_4904;
  wire n_4905, n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912;
  wire n_4913, n_4914, n_4915, n_4916, n_4917, n_4918, n_4919, n_4920;
  wire n_4921, n_4922, n_4923, n_4924, n_4925, n_4926, n_4927, n_4928;
  wire n_4929, n_4930, n_4931, n_4932, n_4933, n_4934, n_4935, n_4936;
  wire n_4937, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944;
  wire n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952;
  wire n_4953, n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960;
  wire n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968;
  wire n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976;
  wire n_4977, n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984;
  wire n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992;
  wire n_4993, n_4994, n_4995, n_4996, n_4997, n_4998, n_4999, n_5000;
  wire n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008;
  wire n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015, n_5016;
  wire n_5017, n_5018, n_5019, n_5020, n_5021, n_5022, n_5023, n_5024;
  wire n_5025, n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032;
  wire n_5033, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040;
  wire n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048;
  wire n_5049, n_5050, n_5051, n_5052, n_5053, n_5054, n_5055, n_5056;
  wire n_5057, n_5058, n_5059, n_5060, n_5061, n_5062, n_5063, n_5064;
  wire n_5065, n_5066, n_5067, n_5068, n_5069, n_5070, n_5071, n_5072;
  wire n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079, n_5080;
  wire n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087, n_5088;
  wire n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095, n_5096;
  wire n_5097, n_5098, n_5099, n_5100, n_5101, n_5102, n_5103, n_5104;
  wire n_5105, n_5106, n_5107, n_5108, n_5109, n_5110, n_5111, n_5112;
  wire n_5113, n_5114, n_5115, n_5116, n_5117, n_5118, n_5119, n_5120;
  wire n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127, n_5128;
  wire n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5136;
  wire n_5137, n_5138, n_5139, n_5140, n_5141, n_5142, n_5143, n_5144;
  wire n_5145, n_5146, n_5147, n_5148, n_5149, n_5150, n_5151, n_5152;
  wire n_5153, n_5154, n_5155, n_5156, n_5157, n_5158, n_5159, n_5160;
  wire n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168;
  wire n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176;
  wire n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5184;
  wire n_5185, n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192;
  wire n_5193, n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200;
  wire n_5201, n_5202, n_5203, n_5204, n_5205, n_5206, n_5207, n_5208;
  wire n_5209, n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5216;
  wire n_5217, n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224;
  wire n_5225, n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232;
  wire n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240;
  wire n_5241, n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, n_5248;
  wire n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256;
  wire n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264;
  wire n_5265, n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272;
  wire n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280;
  wire n_5281, n_5282, n_5283, n_5284, n_5285, n_5286, n_5287, n_5288;
  wire n_5289, n_5290, n_5291, n_5292, n_5293, n_5294, n_5295, n_5296;
  wire n_5297, n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304;
  wire n_5305, n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312;
  wire n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320;
  wire n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328;
  wire n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336;
  wire n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344;
  wire n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352;
  wire n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5360;
  wire n_5361, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367, n_5368;
  wire n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375, n_5376;
  wire n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384;
  wire n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, n_5392;
  wire n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400;
  wire n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408;
  wire n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416;
  wire n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424;
  wire n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432;
  wire n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440;
  wire n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448;
  wire n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456;
  wire n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464;
  wire n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472;
  wire n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480;
  wire n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488;
  wire n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496;
  wire n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504;
  wire n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512;
  wire n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520;
  wire n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528;
  wire n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536;
  wire n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544;
  wire n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552;
  wire n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560;
  wire n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568;
  wire n_5569, n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576;
  wire n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584;
  wire n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592;
  wire n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600;
  wire n_5601, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5627;
  wire n_5628, n_5682, n_5684, n_5686, n_5688, n_5690, n_5692, n_5694;
  wire n_5696, n_5698, n_5700, n_5702, n_5704, n_5705, n_5706, n_5707;
  wire n_5708, n_5709, n_5710, n_5711, n_5712, n_5713, n_5714, n_5715;
  wire n_5716, n_5717, n_5718, n_5719, n_5720, n_5721, n_5722, n_5723;
  wire n_5724, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735;
  wire n_5736, n_5737, n_5738, n_5739, n_5740, n_5741, n_5742, n_5743;
  wire n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, n_5755, n_5756;
  wire n_5757, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764;
  wire n_5765, n_5766, n_5767, n_5768, n_5769, n_5770, n_5771, n_5772;
  wire n_5773, n_5774, n_5775, n_5776, n_5777, n_5778, n_5779, n_5780;
  wire n_5781, n_5782, n_5783, n_5784, n_5785, n_5786, n_5787, n_5788;
  wire n_5789, n_5790, n_5791, n_5792, n_5793, n_5794, n_5795, n_5796;
  wire n_5797, n_5798, n_5799, n_5800, n_5801, n_5802, n_5803, n_5804;
  wire n_5805, n_5806, n_5807, n_5808, n_5809, n_5810, n_5811, n_5812;
  wire n_5813, n_5814, n_5815, n_5816, n_5817, n_5818, n_5819, n_5820;
  wire n_5821, n_5822, n_5823, n_5824, n_5825, n_5826, n_5827, n_5828;
  wire n_5829, n_5830, n_5831, n_5832, n_5833, n_5834, n_5835, n_5836;
  wire n_5837, n_5838, n_5839, n_5840, n_5841, n_5842, n_5843, n_5844;
  wire n_5845, n_5846, n_5847, n_5848, n_5849, n_5850, n_5851, n_5852;
  wire n_5853, n_5854, n_5855, n_5856, n_5857, n_5858, n_5859, n_5860;
  wire n_5861, n_5862, n_5863, n_5864, n_5865, n_5866, n_5867, n_5868;
  wire n_5869, n_5870, n_5871, n_5872, n_5873, n_5874, n_5875, n_5876;
  wire n_5877, n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884;
  wire n_5885, n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892;
  wire n_5893, n_5894, n_5895, n_5896, n_5897, n_5898, n_5899, n_5900;
  wire n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907, n_5908;
  wire n_5909, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915, n_5916;
  wire n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923, n_5924;
  wire n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932;
  wire n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940;
  wire n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5985, n_5987;
  wire n_5988, n_5991, n_5992, n_5993, n_5994, n_5995, n_5996, n_5997;
  wire n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004, n_6005;
  wire n_6006, n_6007, n_6008, n_6010, n_6011, n_6013, n_6014, n_6015;
  wire n_6048, n_6049, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055;
  wire n_6056, n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6063;
  wire n_6064, n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071;
  wire n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079;
  wire n_6080, n_6081, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087;
  wire n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128;
  wire n_6129, n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136;
  wire n_6137, n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144;
  wire n_6145, n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6152;
  wire n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6159, n_6160;
  wire n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167, n_6168;
  wire n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175, n_6176;
  wire n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183, n_6184;
  wire n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192;
  wire n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199, n_6200;
  wire n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207, n_6208;
  wire n_6209, n_6210, n_6211, n_6212, n_6213, n_6214, n_6215, n_6216;
  wire n_6217, n_6218, n_6238, n_6239, n_6240, n_6241, n_6242, n_6243;
  wire n_6244, n_6245, n_6246, n_6247, n_6248, n_6249, n_6250, n_6251;
  wire n_6252, n_6253, n_6254, n_6255, n_6256, n_6257, n_6258, n_6259;
  wire n_6260, n_6261, n_6262, n_6263, n_6264, n_6265, n_6266, n_6267;
  wire n_6268, n_6269, n_6270, n_6271, n_6272, n_6273, n_6274, n_6275;
  wire n_6276, n_6277, n_6278, n_6279, n_6280, n_6281, n_6282, n_6283;
  wire n_6284, n_6285, n_6286, n_6287, n_6288, n_6289, n_6290, n_6291;
  wire n_6292, n_6293, n_6294, n_6295, n_6296, n_6297, n_6298, n_6299;
  wire n_6300, n_6301, n_6302, n_6303, n_6304, n_6305, n_6306, n_6307;
  wire n_6308, n_6309, n_6310, n_6311, n_6312, n_6313, n_6314, n_6315;
  wire n_6316, n_6317, n_6318, n_6319, n_6320, n_6321, n_6322, n_6323;
  wire n_6324, n_6325, n_6326, n_6327, n_6328, n_6329, n_6330, n_6331;
  wire n_6332, n_6333, n_6334, n_6335, n_6336, n_6337, n_6338, n_6339;
  wire n_6340, n_6341, n_6342, n_6343, n_6344, n_6345, n_6346, n_6347;
  wire n_6348, n_6349, n_6350, n_6351, n_6352, n_6353, n_6354, n_6355;
  wire n_6356, n_6357, n_6358, n_6359, n_6360, n_6361, n_6362, n_6363;
  wire n_6364, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370, n_6371;
  wire n_6372, n_6373, n_6374, n_6375, n_6376, n_6377, n_6378, n_6379;
  wire n_6380, n_6381, n_6382, n_6383, n_6384, n_6385, n_6386, n_6387;
  wire n_6388, n_6389, n_6390, n_6391, n_6392, n_6393, n_6394, n_6395;
  wire n_6396, n_6397, n_6398, n_6399, n_6400, n_6401, n_6402, n_6403;
  wire n_6404, n_6405, n_6406, n_6407, n_6408, n_6409, n_6410, n_6411;
  wire n_6412, n_6413, n_6414, n_6415, n_6416, n_6417, n_6418, n_6419;
  wire n_6420, n_6421, n_6422, n_6423, n_6424, n_6425, n_6426, n_6427;
  wire n_6428, n_6429, n_6430, n_6431, n_6432, n_6433, n_6434, n_6435;
  wire n_6436, n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443;
  wire n_6444, n_6445, n_6446, n_6447, n_6448, n_6449, n_6450, n_6451;
  wire n_6452, n_6453, n_6454, n_6455, n_6456, n_6457, n_6458, n_6459;
  wire n_6460, n_6461, n_6462, n_6463, n_6464, n_6465, n_6466, n_6467;
  wire n_6468, n_6469, n_6470, n_6471, n_6472, n_6473, n_6474, n_6475;
  wire n_6476, n_6477, n_6478, n_6479, n_6480, n_6481, n_6482, n_6483;
  wire n_6484, n_6485, n_6486, n_6487, n_6488, n_6489, n_6490, n_6491;
  wire n_6492, n_6493, n_6494, n_6495, n_6496, n_6497, n_6498, n_6499;
  wire n_6500, n_6501, n_6502, n_6503, n_6504, n_6505, n_6506, n_6507;
  wire n_6508, n_6509, n_6510, n_6511, n_6512, n_6513, n_6514, n_6515;
  wire n_6516, n_6517, n_6519, n_6520, n_6522, n_6523, n_6524, n_6525;
  wire n_6526, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532, n_6533;
  wire n_6534, n_6535, n_6536, n_6537, n_6538, n_6539, n_6540, n_6541;
  wire n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548, n_6549;
  wire n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556, n_6557;
  wire n_6558, n_6559, n_6560, n_6561, n_6562, n_6563, n_6564, n_6565;
  wire n_6566, n_6567, n_6568, n_6569, n_6570, n_6571, n_6572, n_6573;
  wire n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, n_6580, n_6581;
  wire n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6588, n_6589;
  wire n_6590, n_6591, n_6593, n_6594, n_6595, n_6596, n_6597, n_6598;
  wire n_6599, n_6600, n_6601, n_6602, n_6603, n_6604, n_6605, n_6606;
  wire n_6607, n_6608, n_6609, n_6610, n_6611, n_6612, n_6613, n_6614;
  wire n_6615, n_6616, n_6617, n_6618, n_6619, n_6620, n_6621, n_6622;
  wire n_6623, n_6624, n_6625, n_6627, n_6628, n_6629, n_6630, n_6631;
  wire n_6632, n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640;
  wire n_6641, n_6642, n_6643, n_6644, n_6645, n_6646, n_6647, n_6648;
  wire n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655, n_6656;
  wire n_6657, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663, n_6664;
  wire n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671, n_6672;
  wire n_6673, n_6674, n_6675, n_6676, n_6677, n_6678, n_6679, n_6680;
  wire n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687, n_6688;
  wire n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695, n_6696;
  wire n_6697, n_6698, n_6699, n_6700, n_6701, n_6702, n_6703, n_6704;
  wire n_6705, n_6706, n_6707, n_6708, n_6710, n_6711, n_6712, n_6713;
  wire n_6714, n_6715, n_6716, n_6717, n_6718, n_6719, n_6720, n_6721;
  wire n_6722, n_6723, n_6724, n_6725, n_6726, n_6729, n_6730, n_6731;
  wire n_6733, n_6734, n_6735, n_6736, n_6737, n_6738, n_6739, n_6740;
  wire n_6741, n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748;
  wire n_6749, n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756;
  wire n_6757, n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764;
  wire n_6765, n_6766, n_6767, n_6768, n_6776, n_6777, n_6778, n_6779;
  wire n_6780, n_6781, n_6782, n_6783, n_6784, n_6785, n_6786, n_6787;
  wire prev_load_request, rc_gclk, rc_gclk_205490, rc_gclk_205493,
       rc_gclk_205496, rc_gclk_205499, rc_gclk_205502, rc_gclk_205505;
  wire rc_gclk_205508, rc_gclk_205511, rc_gclk_205514, rc_gclk_205517,
       rc_gclk_205520, rc_gclk_205523, rc_gclk_205526, rc_gclk_205529;
  wire rc_gclk_205532, rc_gclk_205535, rc_gclk_205538, rc_gclk_205541,
       rc_gclk_205544, rc_gclk_205547, rc_gclk_205550, rc_gclk_205553;
  wire rc_gclk_205556, rc_gclk_205559, rc_gclk_205562, rc_gclk_205565,
       rc_gclk_205568, rc_gclk_205571, rc_gclk_205574, rc_gclk_205577;
  wire rc_gclk_205580, rc_gclk_205583, rc_gclk_205586, rc_gclk_205589,
       rc_gclk_205592, rc_gclk_205595, rc_gclk_205598, rc_gclk_205601;
  wire rc_gclk_205603, rc_gclk_205606, rc_gclk_205610, reset_reg,
       \rs1_data[0]_39306 , \rs1_data[7]_39386 , \rs1_data[8]_39396 ,
       \rs1_data[14]_39466 ;
  wire \rs1_data[15]_39476 , \rs1_data[16]_39486 , \rs1_data[17]_39496
       , \rs1_data[21]_39536 , \rs1_data[22]_39546 ,
       \rs1_data[23]_39246 , \rs1_data[24]_39256 , \rs1_data[26]_39276 ;
  wire \rs1_data[27]_39286 , \rs1_data[28]_39296 , \rs1_data[29]_39336
       , \rs1_data[30]_39446 , store_commit_cycle, store_type,
       system_type, take_trap_39145;
  RC_CG_MOD_AUTO_rvsteel_core RC_CG_HIER_INST1(.ck_in (clock), .enable
       (n_6502), .test (1'b0), .ck_out (rc_gclk));
  RC_CG_MOD_AUTO_rvsteel_core_9 RC_CG_HIER_INST10(.ck_in (clock),
       .enable (n_6493), .test (1'b0), .ck_out (rc_gclk_205514));
  RC_CG_MOD_AUTO_rvsteel_core_10 RC_CG_HIER_INST11(.ck_in (clock),
       .enable (n_6492), .test (1'b0), .ck_out (rc_gclk_205517));
  RC_CG_MOD_AUTO_rvsteel_core_11 RC_CG_HIER_INST12(.ck_in (clock),
       .enable (n_6491), .test (1'b0), .ck_out (rc_gclk_205520));
  RC_CG_MOD_AUTO_rvsteel_core_12 RC_CG_HIER_INST13(.ck_in (clock),
       .enable (n_6490), .test (1'b0), .ck_out (rc_gclk_205523));
  RC_CG_MOD_AUTO_rvsteel_core_13 RC_CG_HIER_INST14(.ck_in (clock),
       .enable (n_6489), .test (1'b0), .ck_out (rc_gclk_205526));
  RC_CG_MOD_AUTO_rvsteel_core_14 RC_CG_HIER_INST15(.ck_in (clock),
       .enable (n_6488), .test (1'b0), .ck_out (rc_gclk_205529));
  RC_CG_MOD_AUTO_rvsteel_core_15 RC_CG_HIER_INST16(.ck_in (clock),
       .enable (n_6487), .test (1'b0), .ck_out (rc_gclk_205532));
  RC_CG_MOD_AUTO_rvsteel_core_16 RC_CG_HIER_INST17(.ck_in (clock),
       .enable (n_6486), .test (1'b0), .ck_out (rc_gclk_205535));
  RC_CG_MOD_AUTO_rvsteel_core_17 RC_CG_HIER_INST18(.ck_in (clock),
       .enable (n_6485), .test (1'b0), .ck_out (rc_gclk_205538));
  RC_CG_MOD_AUTO_rvsteel_core_18 RC_CG_HIER_INST19(.ck_in (clock),
       .enable (n_6484), .test (1'b0), .ck_out (rc_gclk_205541));
  RC_CG_MOD_AUTO_rvsteel_core_1 RC_CG_HIER_INST2(.ck_in (clock),
       .enable (n_6501), .test (1'b0), .ck_out (rc_gclk_205490));
  RC_CG_MOD_AUTO_rvsteel_core_19 RC_CG_HIER_INST20(.ck_in (clock),
       .enable (n_6483), .test (1'b0), .ck_out (rc_gclk_205544));
  RC_CG_MOD_AUTO_rvsteel_core_20 RC_CG_HIER_INST21(.ck_in (clock),
       .enable (n_6482), .test (1'b0), .ck_out (rc_gclk_205547));
  RC_CG_MOD_AUTO_rvsteel_core_21 RC_CG_HIER_INST22(.ck_in (clock),
       .enable (n_6481), .test (1'b0), .ck_out (rc_gclk_205550));
  RC_CG_MOD_AUTO_rvsteel_core_22 RC_CG_HIER_INST23(.ck_in (clock),
       .enable (n_6480), .test (1'b0), .ck_out (rc_gclk_205553));
  RC_CG_MOD_AUTO_rvsteel_core_23 RC_CG_HIER_INST24(.ck_in (clock),
       .enable (n_6479), .test (1'b0), .ck_out (rc_gclk_205556));
  RC_CG_MOD_AUTO_rvsteel_core_24 RC_CG_HIER_INST25(.ck_in (clock),
       .enable (n_6478), .test (1'b0), .ck_out (rc_gclk_205559));
  RC_CG_MOD_AUTO_rvsteel_core_25 RC_CG_HIER_INST26(.ck_in (clock),
       .enable (n_6477), .test (1'b0), .ck_out (rc_gclk_205562));
  RC_CG_MOD_AUTO_rvsteel_core_26 RC_CG_HIER_INST27(.ck_in (clock),
       .enable (n_6476), .test (1'b0), .ck_out (rc_gclk_205565));
  RC_CG_MOD_AUTO_rvsteel_core_27 RC_CG_HIER_INST28(.ck_in (clock),
       .enable (n_6475), .test (1'b0), .ck_out (rc_gclk_205568));
  RC_CG_MOD_AUTO_rvsteel_core_28 RC_CG_HIER_INST29(.ck_in (clock),
       .enable (n_6474), .test (1'b0), .ck_out (rc_gclk_205571));
  RC_CG_MOD_AUTO_rvsteel_core_2 RC_CG_HIER_INST3(.ck_in (clock),
       .enable (n_6500), .test (1'b0), .ck_out (rc_gclk_205493));
  RC_CG_MOD_AUTO_rvsteel_core_29 RC_CG_HIER_INST30(.ck_in (clock),
       .enable (n_6473), .test (1'b0), .ck_out (rc_gclk_205574));
  RC_CG_MOD_AUTO_rvsteel_core_30 RC_CG_HIER_INST31(.ck_in (clock),
       .enable (n_6472), .test (1'b0), .ck_out (rc_gclk_205577));
  RC_CG_MOD_AUTO_rvsteel_core_31 RC_CG_HIER_INST32(.ck_in (clock),
       .enable (n_6471), .test (1'b0), .ck_out (rc_gclk_205580));
  RC_CG_MOD_AUTO_rvsteel_core_32 RC_CG_HIER_INST33(.ck_in (clock),
       .enable (n_6470), .test (1'b0), .ck_out (rc_gclk_205583));
  RC_CG_MOD_AUTO_rvsteel_core_33 RC_CG_HIER_INST34(.ck_in (clock),
       .enable (n_6469), .test (1'b0), .ck_out (rc_gclk_205586));
  RC_CG_MOD_AUTO_rvsteel_core_34 RC_CG_HIER_INST35(.ck_in (clock),
       .enable (n_6468), .test (1'b0), .ck_out (rc_gclk_205589));
  RC_CG_MOD_AUTO_rvsteel_core_35 RC_CG_HIER_INST36(.ck_in (clock),
       .enable (n_6467), .test (1'b0), .ck_out (rc_gclk_205592));
  RC_CG_MOD_AUTO_rvsteel_core_36 RC_CG_HIER_INST37(.ck_in (clock),
       .enable (n_6466), .test (1'b0), .ck_out (rc_gclk_205595));
  RC_CG_MOD_AUTO_rvsteel_core_37 RC_CG_HIER_INST38(.ck_in (clock),
       .enable (n_6465), .test (1'b0), .ck_out (rc_gclk_205598));
  RC_CG_MOD_AUTO_rvsteel_core_38 RC_CG_HIER_INST39(.ck_in (clock),
       .enable (n_6464), .test (1'b0), .ck_out (rc_gclk_205601));
  RC_CG_MOD_AUTO_rvsteel_core_3 RC_CG_HIER_INST4(.ck_in (clock),
       .enable (n_6499), .test (1'b0), .ck_out (rc_gclk_205496));
  RC_CG_MOD_AUTO_rvsteel_core_39 RC_CG_HIER_INST40(.ck_in (clock),
       .enable (n_5628), .test (1'b0), .ck_out (rc_gclk_205603));
  RC_CG_MOD_AUTO_rvsteel_core_40 RC_CG_HIER_INST41(.ck_in (clock),
       .enable (n_6463), .test (1'b0), .ck_out (rc_gclk_205606));
  RC_CG_MOD_AUTO_rvsteel_core_41 RC_CG_HIER_INST42(.ck_in (clock),
       .enable (n_6462), .test (1'b0), .ck_out (rc_gclk_205610));
  RC_CG_MOD_AUTO_rvsteel_core_4 RC_CG_HIER_INST5(.ck_in (clock),
       .enable (n_6498), .test (1'b0), .ck_out (rc_gclk_205499));
  RC_CG_MOD_AUTO_rvsteel_core_5 RC_CG_HIER_INST6(.ck_in (clock),
       .enable (n_6497), .test (1'b0), .ck_out (rc_gclk_205502));
  RC_CG_MOD_AUTO_rvsteel_core_6 RC_CG_HIER_INST7(.ck_in (clock),
       .enable (n_6496), .test (1'b0), .ck_out (rc_gclk_205505));
  RC_CG_MOD_AUTO_rvsteel_core_7 RC_CG_HIER_INST8(.ck_in (clock),
       .enable (n_6495), .test (1'b0), .ck_out (rc_gclk_205508));
  RC_CG_MOD_AUTO_rvsteel_core_8 RC_CG_HIER_INST9(.ck_in (clock),
       .enable (n_6494), .test (1'b0), .ck_out (rc_gclk_205511));
  csa_tree_add_1660_20_group_293 csa_tree_add_1660_20_groupi(.in_0
       ({alu_sra_result[31], n_4485, \rs1_data[29]_39336 ,
       \rs1_data[28]_39296 , \rs1_data[27]_39286 , \rs1_data[26]_39276
       , n_4481, n_4483, \rs1_data[23]_39246 , n_4463, n_4479, n_4486,
       n_4477, n_4478, n_4482, n_4484, \rs1_data[15]_39476 ,
       \rs1_data[14]_39466 , n_4476, n_4475, n_4474, n_4480, n_4487,
       n_4464, n_4460, n_4466, n_4461, n_4465, n_6757, n_6628, n_6629,
       \rs1_data[0]_39306 }), .in_1 ({UNCONNECTED_HIER_Z0,
       UNCONNECTED_HIER_Z, n_6563, n_6564, n_6565, n_6566, n_6567,
       n_6568, n_6569, n_6570, n_6571, n_6572, n_6573, n_6574, n_6575,
       n_6576, n_6577, n_6578, n_6579, n_6580, n_6581, n_6582, n_6583,
       n_6584, n_6585, n_6586, n_6587, n_6588, n_6589, n_6590, n_6591,
       n_6607, n_6593, n_6594}), .in_2 ({UNCONNECTED_HIER_Z33,
       UNCONNECTED_HIER_Z32, UNCONNECTED_HIER_Z31,
       UNCONNECTED_HIER_Z30, UNCONNECTED_HIER_Z29,
       UNCONNECTED_HIER_Z28, UNCONNECTED_HIER_Z27,
       UNCONNECTED_HIER_Z26, UNCONNECTED_HIER_Z25,
       UNCONNECTED_HIER_Z24, UNCONNECTED_HIER_Z23,
       UNCONNECTED_HIER_Z22, UNCONNECTED_HIER_Z21,
       UNCONNECTED_HIER_Z20, UNCONNECTED_HIER_Z19,
       UNCONNECTED_HIER_Z18, UNCONNECTED_HIER_Z17,
       UNCONNECTED_HIER_Z16, UNCONNECTED_HIER_Z15,
       UNCONNECTED_HIER_Z14, UNCONNECTED_HIER_Z13,
       UNCONNECTED_HIER_Z12, UNCONNECTED_HIER_Z11,
       UNCONNECTED_HIER_Z10, UNCONNECTED_HIER_Z9, UNCONNECTED_HIER_Z8,
       UNCONNECTED_HIER_Z7, UNCONNECTED_HIER_Z6, UNCONNECTED_HIER_Z5,
       UNCONNECTED_HIER_Z4, UNCONNECTED_HIER_Z3, UNCONNECTED_HIER_Z2,
       UNCONNECTED_HIER_Z1, alu_operation_code_39061}), .out_0
       ({n_6052, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058,
       n_6059, n_6060, n_6061, n_6062, n_6063, n_6066, n_6068, n_6069,
       n_6070, n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078,
       n_6079, n_6080, n_6081, n_6082, n_6083, n_6084, n_6085, n_6086,
       n_6087}));
  INX1 g28312(.A (alu_2nd_operand[0]), .Q (n_4533));
  INX1 g28313(.A (n_6562), .Q (n_4532));
  BUX1 g28355(.A (\rs1_data[30]_39446 ), .Q (n_4485));
  BUX1 g28373(.A (\rs1_data[16]_39486 ), .Q (n_4484));
  BUX1 g28341(.A (\rs1_data[24]_39256 ), .Q (n_4483));
  BUX1 g28386(.A (\rs1_data[17]_39496 ), .Q (n_4482));
  BUX1 g28344(.A (\rs1_data[21]_39536 ), .Q (n_4479));
  BUX1 g28380(.A (n_6627), .Q (n_4465));
  BUX1 g28334(.A (\rs1_data[22]_39546 ), .Q (n_4463));
  BUX1 g28367(.A (\rs1_data[7]_39386 ), .Q (n_4460));
  BUX1 g28376(.A (\rs1_data[8]_39396 ), .Q (n_4464));
  BUX1 g28402(.A (current_state[2]), .Q (n_4457));
  BUX1 g28403(.A (current_state[3]), .Q (n_4456));
  NA2X1 g40514(.A (n_4441), .B (n_4449), .Q (\rs1_data[22]_39546 ));
  NA2X1 g40515(.A (n_3350), .B (n_3351), .Q (\rs1_data[30]_39446 ));
  NA2X1 g40516(.A (n_3339), .B (n_3336), .Q (n_4486));
  NA2X2 g40517(.A (n_3335), .B (n_3334), .Q (n_4480));
  NA2X1 g40518(.A (n_6630), .B (n_4451), .Q (\rs1_data[29]_39336 ));
  NA2X1 g40519(.A (n_3343), .B (n_3344), .Q (\rs1_data[17]_39496 ));
  NA2X1 g40520(.A (n_3345), .B (n_3342), .Q (\rs1_data[16]_39486 ));
  NA2X2 g40521(.A (n_4454), .B (n_4455), .Q (\rs1_data[28]_39296 ));
  NA2X1 g40522(.A (n_3348), .B (n_3347), .Q (\rs1_data[24]_39256 ));
  NA2X1 g40523(.A (n_6631), .B (n_4450), .Q (alu_sra_result[31]));
  NA2X2 g40524(.A (n_3341), .B (n_3333), .Q (n_4478));
  NA2X1 g40525(.A (n_3340), .B (n_3338), .Q (\rs1_data[21]_39536 ));
  NA2X1 g40526(.A (n_3346), .B (n_3337), .Q (n_4481));
  NA2X2 g40527(.A (n_4437), .B (n_4447), .Q (n_4476));
  NA2X2 g40528(.A (n_4440), .B (n_4444), .Q (n_4487));
  NA2X1 g40529(.A (n_3349), .B (n_3352), .Q (n_4474));
  NA2X2 g40531(.A (n_3331), .B (n_3332), .Q (n_4477));
  NA3X2 g40533(.A (n_4443), .B (n_4411), .C (n_4360), .Q
       (\rs1_data[14]_39466 ));
  NA3X2 g40534(.A (n_4442), .B (n_4390), .C (n_4393), .Q (n_4475));
  NA3X1 g40535(.A (n_4445), .B (n_4417), .C (n_4392), .Q
       (\rs1_data[7]_39386 ));
  NA3X1 g40536(.A (n_4448), .B (n_4416), .C (n_4419), .Q
       (\rs1_data[15]_39476 ));
  NA2X2 g40537(.A (n_4436), .B (n_4432), .Q (\rs1_data[23]_39246 ));
  NA2X1 g40538(.A (n_4446), .B (n_4429), .Q (\rs1_data[27]_39286 ));
  NA2X2 g40539(.A (n_4435), .B (n_4430), .Q (n_4461));
  NA2X1 g40540(.A (n_4433), .B (n_4431), .Q (\rs1_data[26]_39276 ));
  NA2X1 g40542(.A (n_6632), .B (n_4425), .Q (\rs1_data[8]_39396 ));
  NA2X4 g40544(.A (n_6758), .B (n_4420), .Q (\rs1_data[0]_39306 ));
  NA2X1 g40545(.A (n_4439), .B (n_4434), .Q (n_4466));
  AND5X1 g40546(.A (n_6648), .B (n_6661), .C (n_4260), .D (n_4045), .E
       (n_4057), .Q (n_4455));
  AND6X2 g40562(.A (n_4343), .B (n_4167), .C (n_6662), .D (n_4121), .E
       (n_4041), .F (n_4053), .Q (n_4454));
  AND5X1 g40569(.A (n_6653), .B (n_3329), .C (n_4251), .D (n_3994), .E
       (n_3995), .Q (n_4450));
  NO2X1 g40572(.A (n_4418), .B (n_4396), .Q (n_4449));
  NO2X1 g40573(.A (n_4403), .B (n_4406), .Q (n_4448));
  NO2X1 g40574(.A (n_4414), .B (n_4400), .Q (n_4447));
  NO2X1 g40575(.A (n_4386), .B (n_4381), .Q (n_4446));
  NO2X1 g40576(.A (n_6635), .B (n_6634), .Q (n_4445));
  NO2X1 g40577(.A (n_4413), .B (n_4404), .Q (n_4444));
  NO2X1 g40579(.A (n_4401), .B (n_4402), .Q (n_4443));
  NO2X1 g40580(.A (n_4399), .B (n_4410), .Q (n_4442));
  NO3X1 g40581(.A (n_4398), .B (n_4310), .C (n_6698), .Q (n_4441));
  NO3X1 g40582(.A (n_4397), .B (n_4311), .C (n_6699), .Q (n_4440));
  AND5X1 g40583(.A (n_6665), .B (n_3317), .C (n_4244), .D (n_3912), .E
       (n_3952), .Q (n_4439));
  NO2X1 g40586(.A (n_4388), .B (n_4405), .Q (n_4437));
  NO2X1 g40587(.A (n_4387), .B (n_4383), .Q (n_4436));
  NO2X1 g40588(.A (n_4384), .B (n_4382), .Q (n_4435));
  NO2X1 g40589(.A (n_4412), .B (n_6637), .Q (n_4434));
  NO2X1 g40590(.A (n_4385), .B (n_4380), .Q (n_4433));
  NO2X1 g40591(.A (n_4378), .B (n_4379), .Q (n_4432));
  NO2X1 g40592(.A (n_6639), .B (n_6638), .Q (n_4431));
  AND3X1 g40593(.A (n_4377), .B (n_4235), .C (n_4234), .Q (n_4430));
  NO2X1 g40594(.A (n_6640), .B (n_4376), .Q (n_4429));
  NO3X2 g40597(.A (n_4371), .B (n_4249), .C (n_4241), .Q (n_4426));
  NO2X1 g40598(.A (n_6641), .B (n_4372), .Q (n_4425));
  NO3X2 g40601(.A (n_4362), .B (n_4218), .C (n_4208), .Q (n_4422));
  NO3X2 g40603(.A (n_4389), .B (n_4215), .C (n_4209), .Q (n_4420));
  NO2X1 g40604(.A (n_4303), .B (n_3315), .Q (n_4419));
  NA3X1 g40605(.A (n_6664), .B (n_4071), .C (n_4026), .Q (n_4418));
  NO2X1 g40606(.A (n_4307), .B (n_4322), .Q (n_4417));
  NO2X1 g40607(.A (n_4302), .B (n_4320), .Q (n_4416));
  NO2X1 g40608(.A (n_4304), .B (n_4321), .Q (n_4415));
  NA3X1 g40609(.A (n_4330), .B (n_4036), .C (n_4035), .Q (n_4414));
  NA2X1 g40610(.A (n_6779), .B (n_6663), .Q (n_4413));
  NA2X1 g40611(.A (n_4326), .B (n_6666), .Q (n_4412));
  NO2X1 g40612(.A (n_4324), .B (n_4300), .Q (n_4411));
  NA2X1 g40613(.A (n_6672), .B (n_6673), .Q (n_4410));
  NA2X1 g40617(.A (n_6780), .B (n_6680), .Q (n_4406));
  NA2X1 g40618(.A (n_6683), .B (n_6682), .Q (n_4405));
  NA2X1 g40619(.A (n_6667), .B (n_6676), .Q (n_4404));
  NA2X1 g40620(.A (n_3322), .B (n_6642), .Q (n_4403));
  NA2X1 g40621(.A (n_6668), .B (n_6714), .Q (n_4402));
  NA2X1 g40622(.A (n_6669), .B (n_6681), .Q (n_4401));
  NA2X1 g40623(.A (n_6670), .B (n_6684), .Q (n_4400));
  NA3X1 g40624(.A (n_6671), .B (n_3929), .C (n_3969), .Q (n_4399));
  NA2X1 g40625(.A (n_6675), .B (n_6685), .Q (n_4398));
  NA2X1 g40626(.A (n_6674), .B (n_6686), .Q (n_4397));
  NA2X1 g40627(.A (n_6677), .B (n_6687), .Q (n_4396));
  NO2X1 g40630(.A (n_4313), .B (n_4248), .Q (n_4393));
  AND3X1 g40631(.A (n_4070), .B (n_4023), .C (n_4245), .Q (n_4392));
  AND3X1 g40632(.A (n_4066), .B (n_4014), .C (n_4243), .Q (n_4391));
  NO2X1 g40633(.A (n_4312), .B (n_4323), .Q (n_4390));
  NA3X1 g40634(.A (n_4279), .B (n_3765), .C (n_3778), .Q (n_4389));
  NA3X1 g40635(.A (n_4061), .B (n_4004), .C (n_4239), .Q (n_4388));
  NA2X1 g40636(.A (n_6690), .B (n_6693), .Q (n_4387));
  NA2X1 g40637(.A (n_6694), .B (n_6691), .Q (n_4386));
  NA2X1 g40638(.A (n_6695), .B (n_6692), .Q (n_4385));
  NA3X1 g40639(.A (n_6696), .B (n_3882), .C (n_3883), .Q (n_4384));
  NA3X1 g40640(.A (n_3891), .B (n_3890), .C (n_6759), .Q (n_4383));
  NA3X1 g40641(.A (n_3884), .B (n_3885), .C (n_6782), .Q (n_4382));
  NA3X1 g40642(.A (n_3878), .B (n_3877), .C (n_6783), .Q (n_4381));
  NA3X1 g40643(.A (n_3871), .B (n_3872), .C (n_6710), .Q (n_4380));
  NA2X1 g40644(.A (n_6700), .B (n_6704), .Q (n_4379));
  NA2X1 g40645(.A (n_6701), .B (n_6705), .Q (n_4378));
  NO2X1 g40646(.A (n_4236), .B (n_6706), .Q (n_4377));
  NA2X1 g40647(.A (n_6702), .B (n_6707), .Q (n_4376));
  NA3X1 g40651(.A (n_6784), .B (n_3818), .C (n_3812), .Q (n_4372));
  NA3X2 g40652(.A (n_4200), .B (n_3815), .C (n_3808), .Q (n_4371));
  NO2X1 g40656(.A (n_4217), .B (n_4207), .Q (n_4367));
  NO2X1 g40657(.A (n_4204), .B (n_4213), .Q (n_4366));
  NA3X2 g40661(.A (n_4199), .B (n_3772), .C (n_3781), .Q (n_4362));
  NA3X1 g40662(.A (n_4198), .B (n_3768), .C (n_3777), .Q (n_4361));
  NO2X1 g40663(.A (n_4301), .B (n_4240), .Q (n_4360));
  AN221X1 g40665(.A (n_5113), .B (n_3510), .C (n_5112), .D (n_3526), .E
       (n_4177), .Q (n_4358));
  AN221X1 g40667(.A (n_5435), .B (n_3553), .C (n_5436), .D (n_3554), .E
       (n_4186), .Q (n_4356));
  AN221X1 g40668(.A (n_5445), .B (n_3536), .C (n_5446), .D (n_3546), .E
       (n_4185), .Q (n_4355));
  AN221X1 g40671(.A (n_5109), .B (n_3301), .C (n_5110), .D (n_3512), .E
       (n_4178), .Q (n_4352));
  AND2X1 g40679(.A (n_4126), .B (n_4125), .Q (n_4344));
  AND2X2 g40680(.A (n_4123), .B (n_4122), .Q (n_4343));
  AN221X1 g40685(.A (n_5125), .B (n_3553), .C (n_5126), .D (n_3554), .E
       (n_4139), .Q (n_4338));
  NO2X1 g40690(.A (n_4088), .B (n_4094), .Q (n_4333));
  AND2X1 g40692(.A (n_4143), .B (n_4144), .Q (n_4331));
  NO2X1 g40693(.A (n_4034), .B (n_4075), .Q (n_4330));
  AND2X1 g40694(.A (n_4087), .B (n_4116), .Q (n_4329));
  AND2X1 g40695(.A (n_4113), .B (n_4114), .Q (n_4328));
  NO2X1 g40697(.A (n_4015), .B (n_4067), .Q (n_4326));
  OR4X1 g40699(.A (n_3663), .B (n_3664), .C (n_3665), .D (n_3666), .Q
       (n_4324));
  OR4X1 g40700(.A (n_3689), .B (n_3691), .C (n_3690), .D (n_3710), .Q
       (n_4323));
  NA2X1 g40701(.A (n_4069), .B (n_4022), .Q (n_4322));
  NA2X1 g40702(.A (n_4012), .B (n_4013), .Q (n_4321));
  OR4X1 g40703(.A (n_3675), .B (n_3677), .C (n_3676), .D (n_3702), .Q
       (n_4320));
  AND2X1 g40706(.A (n_4043), .B (n_4044), .Q (n_4317));
  AND2X1 g40708(.A (n_4038), .B (n_4050), .Q (n_4315));
  AND2X1 g40709(.A (n_4040), .B (n_4052), .Q (n_4314));
  OR4X1 g40717(.A (n_3711), .B (n_3712), .C (n_3713), .D (n_3714), .Q
       (n_4313));
  OR4X1 g40718(.A (n_3688), .B (n_3686), .C (n_3687), .D (n_3283), .Q
       (n_4312));
  NA2X1 g40719(.A (n_4074), .B (n_4030), .Q (n_4311));
  NA2X1 g40720(.A (n_4073), .B (n_4032), .Q (n_4310));
  NA2X1 g40723(.A (n_4020), .B (n_4021), .Q (n_4307));
  NA2X1 g40726(.A (n_4065), .B (n_4011), .Q (n_4304));
  NA2X1 g40727(.A (n_4062), .B (n_4005), .Q (n_4303));
  OR4X1 g40728(.A (n_3673), .B (n_3671), .C (n_3672), .D (n_3674), .Q
       (n_4302));
  OR4X1 g40729(.A (n_3696), .B (n_3698), .C (n_3697), .D (n_3699), .Q
       (n_4301));
  OR4X1 g40730(.A (n_3667), .B (n_3668), .C (n_3669), .D (n_3695), .Q
       (n_4300));
  AND2X1 g40752(.A (n_3904), .B (n_3944), .Q (n_4284));
  AND2X1 g40753(.A (n_3902), .B (n_3903), .Q (n_4283));
  AN221X1 g40756(.A (n_5432), .B (n_3295), .C (n_5418), .D (n_3505), .E
       (n_4187), .Q (n_4280));
  NO3X1 g40757(.A (n_3559), .B (n_3558), .C (n_3564), .Q (n_4279));
  AN222X1 g40761(.A (n_3524), .B (n_5425), .C (n_5426), .D (n_3514), .E
       (n_5421), .F (n_3520), .Q (n_4275));
  AN222X1 g40769(.A (n_3518), .B (n_5117), .C (n_5118), .D (n_3517), .E
       (n_5111), .F (n_3520), .Q (n_4268));
  AN222X1 g40770(.A (n_3518), .B (n_5179), .C (n_5180), .D (n_3517), .E
       (n_5173), .F (n_3520), .Q (n_4267));
  AN221X1 g40771(.A (n_5328), .B (n_3520), .C (n_5334), .D (n_3518), .E
       (n_3758), .Q (n_4266));
  AN221X1 g40772(.A (n_5297), .B (n_3520), .C (n_5303), .D (n_3518), .E
       (n_3755), .Q (n_4265));
  AN221X1 g40773(.A (n_4584), .B (n_3520), .C (n_4590), .D (n_3518), .E
       (n_3754), .Q (n_4264));
  AN211X1 g40777(.A (n_3520), .B (n_4708), .C (n_3749), .D (n_3750), .Q
       (n_4260));
  AN221X1 g40778(.A (n_5452), .B (n_3520), .C (n_5458), .D (n_3518), .E
       (n_3747), .Q (n_4259));
  AN221X1 g40779(.A (n_4615), .B (n_3520), .C (n_4621), .D (n_3518), .E
       (n_3745), .Q (n_4258));
  AN211X1 g40784(.A (n_3520), .B (n_4832), .C (n_3735), .D (n_3736), .Q
       (n_4253));
  AN211X1 g40786(.A (n_3520), .B (n_5514), .C (n_3727), .D (n_3728), .Q
       (n_4251));
  AN221X1 g40787(.A (n_5359), .B (n_3520), .C (n_5365), .D (n_3518), .E
       (n_3724), .Q (n_4250));
  NA2X1 g40788(.A (n_3806), .B (n_3813), .Q (n_4249));
  NA3X1 g40789(.A (n_3715), .B (n_3716), .C (n_3692), .Q (n_4248));
  AN211X1 g40793(.A (n_3520), .B (n_4987), .C (n_3708), .D (n_3709), .Q
       (n_4245));
  NO2X1 g40794(.A (n_4019), .B (n_3678), .Q (n_4244));
  AN211X1 g40795(.A (n_3520), .B (n_4894), .C (n_3705), .D (n_3704), .Q
       (n_4243));
  AN21X1 g40796(.A (n_3520), .B (n_5390), .C (n_4010), .Q (n_4242));
  NA2X1 g40797(.A (n_3807), .B (n_3814), .Q (n_4241));
  NA3X1 g40799(.A (n_3700), .B (n_3701), .C (n_3670), .Q (n_4240));
  AN211X1 g40800(.A (n_3520), .B (n_5204), .C (n_3693), .D (n_3694), .Q
       (n_4239));
  NA2X1 g40803(.A (n_3861), .B (n_3862), .Q (n_4236));
  AND2X1 g40804(.A (n_3840), .B (n_3860), .Q (n_4235));
  AND2X1 g40805(.A (n_3839), .B (n_3859), .Q (n_4234));
  AND2X1 g40815(.A (n_3843), .B (n_3844), .Q (n_4227));
  NA2X1 g40823(.A (n_3821), .B (n_3822), .Q (n_4223));
  NA2X1 g40828(.A (n_3779), .B (n_3780), .Q (n_4218));
  NA2X1 g40829(.A (n_3776), .B (n_3775), .Q (n_4217));
  NA2X1 g40831(.A (n_3792), .B (n_3793), .Q (n_4215));
  NA2X1 g40833(.A (n_3788), .B (n_3796), .Q (n_4213));
  NA2X1 g40837(.A (n_3782), .B (n_3783), .Q (n_4209));
  NA2X1 g40838(.A (n_3770), .B (n_3771), .Q (n_4208));
  NA2X1 g40839(.A (n_3766), .B (n_3767), .Q (n_4207));
  NA2X1 g40840(.A (n_3979), .B (n_3764), .Q (n_4206));
  NA2X1 g40842(.A (n_3794), .B (n_3795), .Q (n_4204));
  NO2X2 g40843(.A (n_3799), .B (n_3791), .Q (n_4203));
  NA2X1 g40844(.A (n_3786), .B (n_3800), .Q (n_4202));
  NO2X2 g40846(.A (n_3809), .B (n_3589), .Q (n_4200));
  NO3X2 g40847(.A (n_3560), .B (n_3561), .C (n_3562), .Q (n_4199));
  NO2X1 g40848(.A (n_3769), .B (n_3563), .Q (n_4198));
  AN22X1 g40850(.A (n_3549), .B (n_4844), .C (n_3551), .D (n_4845), .Q
       (n_4196));
  AN22X1 g40851(.A (n_3510), .B (n_5423), .C (n_3526), .D (n_5422), .Q
       (n_4195));
  AN22X1 g40852(.A (n_3508), .B (n_5424), .C (n_3305), .D (n_5429), .Q
       (n_4194));
  AO22X1 g40854(.A (n_3510), .B (n_5175), .C (n_3526), .D (n_5174), .Q
       (n_4192));
  AN22X1 g40855(.A (n_3542), .B (n_5437), .C (n_3544), .D (n_5438), .Q
       (n_4191));
  AN22X1 g40856(.A (n_3538), .B (n_5439), .C (n_3540), .D (n_5440), .Q
       (n_4190));
  AN22X1 g40857(.A (n_3547), .B (n_5447), .C (n_3504), .D (n_5448), .Q
       (n_4189));
  AN22X1 g40858(.A (n_3518), .B (n_5427), .C (n_3517), .D (n_5428), .Q
       (n_4188));
  AO22X1 g40859(.A (n_3522), .B (n_5431), .C (n_3298), .D (n_5430), .Q
       (n_4187));
  AO22X1 g40860(.A (n_3549), .B (n_5433), .C (n_3551), .D (n_5434), .Q
       (n_4186));
  AO22X1 g40861(.A (n_6768), .B (n_5443), .C (n_6767), .D (n_5444), .Q
       (n_4185));
  AN22X1 g40862(.A (n_3548), .B (n_5441), .C (n_3557), .D (n_5442), .Q
       (n_4184));
  NA2X1 g40863(.A (n_3761), .B (n_3762), .Q (n_4183));
  AO22X1 g40865(.A (n_3301), .B (n_5295), .C (n_3512), .D (n_5296), .Q
       (n_4181));
  AN22X1 g40867(.A (n_3301), .B (n_4582), .C (n_3512), .D (n_4583), .Q
       (n_4179));
  ON22X1 g40868(.A (n_3525), .B (n_3365), .C (n_3515), .D (n_3357), .Q
       (n_4178));
  ON22X1 g40869(.A (n_3294), .B (n_3380), .C (n_3506), .D (n_3375), .Q
       (n_4177));
  AN22X1 g40870(.A (n_3508), .B (n_5114), .C (n_3305), .D (n_5119), .Q
       (n_4176));
  AN22X1 g40871(.A (n_3522), .B (n_5121), .C (n_3298), .D (n_5120), .Q
       (n_4175));
  AO22X1 g40872(.A (n_3524), .B (n_5177), .C (n_3514), .D (n_5178), .Q
       (n_4174));
  AN22X1 g40874(.A (n_3508), .B (n_5176), .C (n_3305), .D (n_5181), .Q
       (n_4172));
  AN22X1 g40875(.A (n_3522), .B (n_5183), .C (n_3298), .D (n_5182), .Q
       (n_4171));
  NA2X1 g40877(.A (n_3753), .B (n_3752), .Q (n_4169));
  AN22X1 g40878(.A (n_3510), .B (n_5454), .C (n_3526), .D (n_5453), .Q
       (n_4168));
  AN22X1 g40879(.A (n_3510), .B (n_4710), .C (n_3526), .D (n_4709), .Q
       (n_4167));
  AO22X1 g40880(.A (n_3301), .B (n_4613), .C (n_3512), .D (n_4614), .Q
       (n_4166));
  AN22X1 g40881(.A (n_3510), .B (n_4617), .C (n_3508), .D (n_4618), .Q
       (n_4165));
  AO22X1 g40882(.A (n_3295), .B (n_4595), .C (n_3508), .D (n_4587), .Q
       (n_4164));
  AN22X1 g40885(.A (n_3295), .B (n_5339), .C (n_3505), .D (n_5325), .Q
       (n_4161));
  AN22X1 g40886(.A (n_3522), .B (n_5338), .C (n_3298), .D (n_5337), .Q
       (n_4160));
  AO22X1 g40887(.A (n_3509), .B (n_5331), .C (n_3305), .D (n_5336), .Q
       (n_4159));
  AO22X1 g40889(.A (n_3305), .B (n_5305), .C (n_3505), .D (n_5294), .Q
       (n_4157));
  AN22X1 g40890(.A (n_3295), .B (n_5308), .C (n_3526), .D (n_5298), .Q
       (n_4156));
  AN22X1 g40891(.A (n_3522), .B (n_5307), .C (n_3298), .D (n_5306), .Q
       (n_4155));
  AN22X1 g40892(.A (n_3524), .B (n_4588), .C (n_3514), .D (n_4589), .Q
       (n_4154));
  AN22X1 g40893(.A (n_3522), .B (n_4594), .C (n_3505), .D (n_4581), .Q
       (n_4153));
  AN22X1 g40894(.A (n_3510), .B (n_4586), .C (n_3298), .D (n_4593), .Q
       (n_4152));
  AN22X1 g40895(.A (n_3538), .B (n_5191), .C (n_3540), .D (n_5192), .Q
       (n_4151));
  AN22X1 g40896(.A (n_3536), .B (n_5135), .C (n_3546), .D (n_5136), .Q
       (n_4150));
  AN22X1 g40897(.A (n_3547), .B (n_5137), .C (n_3504), .D (n_5138), .Q
       (n_4149));
  AN22X1 g40898(.A (n_3542), .B (n_5127), .C (n_3544), .D (n_5128), .Q
       (n_4148));
  AN22X1 g40899(.A (n_3538), .B (n_5129), .C (n_3540), .D (n_5130), .Q
       (n_4147));
  AN22X1 g40900(.A (n_3536), .B (n_5197), .C (n_3546), .D (n_5198), .Q
       (n_4146));
  AN22X1 g40901(.A (n_3547), .B (n_5199), .C (n_3504), .D (n_5200), .Q
       (n_4145));
  AN22X1 g40902(.A (n_3542), .B (n_5189), .C (n_3544), .D (n_5190), .Q
       (n_4144));
  AN22X1 g40903(.A (n_3553), .B (n_5187), .C (n_3554), .D (n_5188), .Q
       (n_4143));
  AN22X1 g40904(.A (n_3549), .B (n_5185), .C (n_3551), .D (n_5186), .Q
       (n_4142));
  AN22X1 g40905(.A (n_6768), .B (n_5133), .C (n_6767), .D (n_5134), .Q
       (n_4141));
  AN22X1 g40906(.A (n_3548), .B (n_5131), .C (n_3557), .D (n_5132), .Q
       (n_4140));
  AO22X1 g40907(.A (n_3549), .B (n_5123), .C (n_3551), .D (n_5124), .Q
       (n_4139));
  AN22X1 g40908(.A (n_3548), .B (n_5193), .C (n_3557), .D (n_5194), .Q
       (n_4138));
  AN22X1 g40909(.A (n_6768), .B (n_5195), .C (n_6767), .D (n_5196), .Q
       (n_4137));
  AO22X1 g40911(.A (n_3301), .B (n_5078), .C (n_3512), .D (n_5079), .Q
       (n_4135));
  NA2X1 g40913(.A (n_3738), .B (n_3739), .Q (n_4133));
  ON22X1 g40914(.A (n_3300), .B (n_3359), .C (n_3513), .D (n_3353), .Q
       (n_4132));
  AO22X1 g40915(.A (n_3301), .B (n_5357), .C (n_3512), .D (n_5358), .Q
       (n_4131));
  AN22X1 g40916(.A (n_3510), .B (n_5361), .C (n_3526), .D (n_5360), .Q
       (n_4130));
  ON22X1 g40917(.A (n_3511), .B (n_3381), .C (n_3527), .D (n_3369), .Q
       (n_4129));
  ON22X1 g40919(.A (n_3525), .B (n_3355), .C (n_3515), .D (n_3362), .Q
       (n_4127));
  AN22X1 g40920(.A (n_3295), .B (n_5463), .C (n_3505), .D (n_5449), .Q
       (n_4126));
  AN22X1 g40921(.A (n_3522), .B (n_5462), .C (n_3298), .D (n_5461), .Q
       (n_4125));
  AN22X1 g40922(.A (n_3508), .B (n_5455), .C (n_3305), .D (n_5460), .Q
       (n_4124));
  AN21X1 g40923(.A (n_3295), .B (n_4719), .C (n_3751), .Q (n_4123));
  AN21X1 g40924(.A (n_3522), .B (n_4718), .C (n_3744), .Q (n_4122));
  AN22X1 g40925(.A (n_3508), .B (n_4711), .C (n_3305), .D (n_4716), .Q
       (n_4121));
  AN22X1 g40927(.A (n_3305), .B (n_4623), .C (n_3298), .D (n_4624), .Q
       (n_4119));
  AN22X1 g40928(.A (n_3295), .B (n_4626), .C (n_3526), .D (n_4616), .Q
       (n_4118));
  AN22X1 g40929(.A (n_3522), .B (n_4625), .C (n_3505), .D (n_4612), .Q
       (n_4117));
  AN22X1 g40930(.A (n_3549), .B (n_4596), .C (n_3551), .D (n_4597), .Q
       (n_4116));
  AN22X1 g40931(.A (n_3553), .B (n_4598), .C (n_3554), .D (n_4599), .Q
       (n_4115));
  AN22X1 g40932(.A (n_3548), .B (n_4604), .C (n_3557), .D (n_4605), .Q
       (n_4114));
  AN22X1 g40933(.A (n_6768), .B (n_4606), .C (n_6767), .D (n_4607), .Q
       (n_4113));
  AN22X1 g40934(.A (n_6768), .B (n_5350), .C (n_6767), .D (n_5351), .Q
       (n_4112));
  AN22X1 g40935(.A (n_3548), .B (n_5348), .C (n_3557), .D (n_5349), .Q
       (n_4111));
  AO22X1 g40936(.A (n_3553), .B (n_5342), .C (n_3554), .D (n_5343), .Q
       (n_4110));
  AN22X1 g40937(.A (n_3549), .B (n_5340), .C (n_3551), .D (n_5341), .Q
       (n_4109));
  AN22X1 g40938(.A (n_3548), .B (n_5317), .C (n_3557), .D (n_5318), .Q
       (n_4108));
  AN22X1 g40939(.A (n_6768), .B (n_5319), .C (n_6767), .D (n_5320), .Q
       (n_4107));
  AO22X1 g40940(.A (n_3549), .B (n_5309), .C (n_3551), .D (n_5310), .Q
       (n_4106));
  AN22X1 g40941(.A (n_3553), .B (n_5311), .C (n_3554), .D (n_5312), .Q
       (n_4105));
  NA2X1 g40942(.A (n_3734), .B (n_3733), .Q (n_4104));
  NA2X1 g40945(.A (n_3721), .B (n_3743), .Q (n_4101));
  AO22X1 g40947(.A (n_3509), .B (n_5083), .C (n_3305), .D (n_5088), .Q
       (n_4099));
  AO22X1 g40948(.A (n_3522), .B (n_5090), .C (n_3298), .D (n_5089), .Q
       (n_4098));
  NA2X1 g40952(.A (n_3719), .B (n_3737), .Q (n_4094));
  AN22X1 g40954(.A (n_3295), .B (n_5370), .C (n_3505), .D (n_5356), .Q
       (n_4092));
  AN22X1 g40955(.A (n_3522), .B (n_5369), .C (n_3298), .D (n_5368), .Q
       (n_4091));
  AN22X1 g40956(.A (n_3508), .B (n_5362), .C (n_3305), .D (n_5367), .Q
       (n_4090));
  ON22X1 g40958(.A (n_3523), .B (n_3377), .C (n_3297), .D (n_3379), .Q
       (n_4088));
  AN22X1 g40959(.A (n_3542), .B (n_4600), .C (n_3544), .D (n_4601), .Q
       (n_4087));
  AN22X1 g40960(.A (n_3538), .B (n_4602), .C (n_3540), .D (n_4603), .Q
       (n_4086));
  AN22X1 g40961(.A (n_3536), .B (n_4608), .C (n_3546), .D (n_4609), .Q
       (n_4085));
  AN22X1 g40962(.A (n_3547), .B (n_4610), .C (n_3504), .D (n_4611), .Q
       (n_4084));
  AN22X1 g40963(.A (n_3536), .B (n_5352), .C (n_3546), .D (n_5353), .Q
       (n_4083));
  AN22X1 g40964(.A (n_3547), .B (n_5354), .C (n_3504), .D (n_5355), .Q
       (n_4082));
  AN22X1 g40966(.A (n_3538), .B (n_5346), .C (n_3540), .D (n_5347), .Q
       (n_4080));
  AN22X1 g40967(.A (n_3536), .B (n_5321), .C (n_3546), .D (n_5322), .Q
       (n_4079));
  AN22X1 g40968(.A (n_3547), .B (n_5323), .C (n_3504), .D (n_5324), .Q
       (n_4078));
  AN22X1 g40970(.A (n_3538), .B (n_5315), .C (n_3540), .D (n_5316), .Q
       (n_4076));
  AO22X1 g40971(.A (n_3510), .B (n_5206), .C (n_3526), .D (n_5205), .Q
       (n_4075));
  AN22X1 g40972(.A (n_3301), .B (n_5047), .C (n_3512), .D (n_5048), .Q
       (n_4074));
  AN22X1 g40973(.A (n_3301), .B (n_5481), .C (n_3512), .D (n_5482), .Q
       (n_4073));
  ON22X1 g40974(.A (n_3511), .B (n_3376), .C (n_3527), .D (n_3354), .Q
       (n_4072));
  AN22X1 g40975(.A (n_3510), .B (n_5485), .C (n_3526), .D (n_5484), .Q
       (n_4071));
  AN22X1 g40976(.A (n_3301), .B (n_4985), .C (n_3512), .D (n_4986), .Q
       (n_4070));
  AN22X1 g40977(.A (n_3510), .B (n_4989), .C (n_3509), .D (n_4990), .Q
       (n_4069));
  AO22X1 g40979(.A (n_3510), .B (n_4958), .C (n_3526), .D (n_4957), .Q
       (n_4067));
  AN22X1 g40980(.A (n_3301), .B (n_4892), .C (n_3512), .D (n_4893), .Q
       (n_4066));
  AN22X1 g40981(.A (n_3510), .B (n_4896), .C (n_3526), .D (n_4895), .Q
       (n_4065));
  AN22X1 g40982(.A (n_3301), .B (n_5388), .C (n_3512), .D (n_5389), .Q
       (n_4064));
  AN22X1 g40983(.A (n_3510), .B (n_5392), .C (n_3526), .D (n_5391), .Q
       (n_4063));
  AN22X1 g40984(.A (n_3301), .B (n_5264), .C (n_3512), .D (n_5265), .Q
       (n_4062));
  AN22X1 g40985(.A (n_3301), .B (n_5202), .C (n_3512), .D (n_5203), .Q
       (n_4061));
  AN22X1 g40986(.A (n_3542), .B (n_5468), .C (n_3544), .D (n_5469), .Q
       (n_4060));
  AN22X1 g40988(.A (n_3538), .B (n_5470), .C (n_3540), .D (n_5471), .Q
       (n_4058));
  AN22X1 g40989(.A (n_3547), .B (n_4734), .C (n_3504), .D (n_4735), .Q
       (n_4057));
  AN22X1 g40990(.A (n_3536), .B (n_5476), .C (n_3546), .D (n_5477), .Q
       (n_4056));
  AN22X1 g40991(.A (n_3547), .B (n_5478), .C (n_3504), .D (n_5479), .Q
       (n_4055));
  AN22X1 g40993(.A (n_3538), .B (n_4726), .C (n_3540), .D (n_4727), .Q
       (n_4053));
  AN22X1 g40994(.A (n_3542), .B (n_4631), .C (n_3544), .D (n_4632), .Q
       (n_4052));
  AN22X1 g40995(.A (n_3538), .B (n_4633), .C (n_3540), .D (n_4634), .Q
       (n_4051));
  AN22X1 g40996(.A (n_3536), .B (n_4639), .C (n_3546), .D (n_4640), .Q
       (n_4050));
  AN22X1 g40997(.A (n_3547), .B (n_4641), .C (n_3504), .D (n_4642), .Q
       (n_4049));
  AN22X1 g40998(.A (n_3549), .B (n_5464), .C (n_3551), .D (n_5465), .Q
       (n_4048));
  AO22X1 g40999(.A (n_3548), .B (n_4728), .C (n_3557), .D (n_4729), .Q
       (n_4047));
  AN22X1 g41000(.A (n_3553), .B (n_5466), .C (n_3554), .D (n_5467), .Q
       (n_4046));
  AN22X1 g41001(.A (n_6768), .B (n_4730), .C (n_6767), .D (n_4731), .Q
       (n_4045));
  AN22X1 g41002(.A (n_3548), .B (n_5472), .C (n_3557), .D (n_5473), .Q
       (n_4044));
  AN22X1 g41003(.A (n_6768), .B (n_5474), .C (n_6767), .D (n_5475), .Q
       (n_4043));
  AO22X1 g41004(.A (n_3549), .B (n_4720), .C (n_3551), .D (n_4721), .Q
       (n_4042));
  AN22X1 g41005(.A (n_3553), .B (n_4722), .C (n_3554), .D (n_4723), .Q
       (n_4041));
  AN22X1 g41006(.A (n_3553), .B (n_4629), .C (n_3554), .D (n_4630), .Q
       (n_4040));
  AN22X1 g41007(.A (n_3549), .B (n_4627), .C (n_3551), .D (n_4628), .Q
       (n_4039));
  AN22X1 g41008(.A (n_3548), .B (n_4635), .C (n_3557), .D (n_4636), .Q
       (n_4038));
  AN22X1 g41009(.A (n_6768), .B (n_4637), .C (n_6767), .D (n_4638), .Q
       (n_4037));
  AN22X1 g41010(.A (n_3295), .B (n_5215), .C (n_3505), .D (n_5201), .Q
       (n_4036));
  AN22X1 g41011(.A (n_3522), .B (n_5214), .C (n_3298), .D (n_5213), .Q
       (n_4035));
  AO22X1 g41012(.A (n_3509), .B (n_5207), .C (n_3305), .D (n_5212), .Q
       (n_4034));
  AN22X1 g41014(.A (n_3524), .B (n_5487), .C (n_3514), .D (n_5488), .Q
       (n_4032));
  AN22X1 g41016(.A (n_3524), .B (n_5053), .C (n_3514), .D (n_5054), .Q
       (n_4030));
  AO22X1 g41018(.A (n_3522), .B (n_5059), .C (n_3298), .D (n_5058), .Q
       (n_4028));
  AN22X1 g41020(.A (n_3295), .B (n_5494), .C (n_3505), .D (n_5480), .Q
       (n_4026));
  NA2X1 g41021(.A (n_3682), .B (n_3681), .Q (n_4025));
  AN22X1 g41023(.A (n_3524), .B (n_4991), .C (n_3514), .D (n_4992), .Q
       (n_4023));
  AN22X1 g41024(.A (n_3305), .B (n_4995), .C (n_3505), .D (n_4984), .Q
       (n_4022));
  AN22X1 g41025(.A (n_3295), .B (n_4998), .C (n_3298), .D (n_4996), .Q
       (n_4021));
  AN22X1 g41026(.A (n_3522), .B (n_4997), .C (n_3526), .D (n_4988), .Q
       (n_4020));
  ON22X1 g41027(.A (n_3519), .B (n_3364), .C (n_3302), .D (n_3370), .Q
       (n_4019));
  NA2X1 g41028(.A (n_3706), .B (n_3707), .Q (n_4018));
  ON22X1 g41029(.A (n_3294), .B (n_3374), .C (n_3506), .D (n_3373), .Q
       (n_4017));
  AO22X1 g41031(.A (n_3509), .B (n_4959), .C (n_3305), .D (n_4964), .Q
       (n_4015));
  AN22X1 g41032(.A (n_3518), .B (n_4900), .C (n_3517), .D (n_4901), .Q
       (n_4014));
  AN22X1 g41033(.A (n_3296), .B (n_4905), .C (n_3505), .D (n_4891), .Q
       (n_4013));
  AN22X1 g41034(.A (n_3509), .B (n_4897), .C (n_3305), .D (n_4902), .Q
       (n_4012));
  AN22X1 g41035(.A (n_3522), .B (n_4904), .C (n_3298), .D (n_4903), .Q
       (n_4011));
  ON22X1 g41036(.A (n_3519), .B (n_3356), .C (n_3302), .D (n_3358), .Q
       (n_4010));
  AN22X1 g41037(.A (n_3524), .B (n_5394), .C (n_3514), .D (n_5395), .Q
       (n_4009));
  AN22X1 g41038(.A (n_3295), .B (n_5401), .C (n_3505), .D (n_5387), .Q
       (n_4008));
  AN22X1 g41039(.A (n_3509), .B (n_5393), .C (n_3305), .D (n_5398), .Q
       (n_4007));
  AN22X1 g41040(.A (n_3522), .B (n_5400), .C (n_3298), .D (n_5399), .Q
       (n_4006));
  AN22X1 g41041(.A (n_3524), .B (n_5270), .C (n_3514), .D (n_5271), .Q
       (n_4005));
  AN22X1 g41042(.A (n_3524), .B (n_5208), .C (n_3514), .D (n_5209), .Q
       (n_4004));
  AN22X1 g41043(.A (n_3536), .B (n_4856), .C (n_3546), .D (n_4857), .Q
       (n_4003));
  AN22X1 g41044(.A (n_3547), .B (n_4858), .C (n_3504), .D (n_4859), .Q
       (n_4002));
  AN22X1 g41045(.A (n_3536), .B (n_5104), .C (n_3546), .D (n_5105), .Q
       (n_4001));
  AN22X1 g41046(.A (n_3547), .B (n_5106), .C (n_3504), .D (n_5107), .Q
       (n_4000));
  AN22X1 g41047(.A (n_3542), .B (n_5096), .C (n_3544), .D (n_5097), .Q
       (n_3999));
  AN22X1 g41048(.A (n_3538), .B (n_5098), .C (n_3540), .D (n_5099), .Q
       (n_3998));
  AN22X1 g41049(.A (n_3542), .B (n_4848), .C (n_3544), .D (n_4849), .Q
       (n_3997));
  AN22X1 g41050(.A (n_3538), .B (n_4850), .C (n_3540), .D (n_4851), .Q
       (n_3996));
  AN22X1 g41051(.A (n_3536), .B (n_5538), .C (n_3546), .D (n_5539), .Q
       (n_3995));
  AN22X1 g41052(.A (n_3547), .B (n_5540), .C (n_3504), .D (n_5541), .Q
       (n_3994));
  AN22X1 g41053(.A (n_3542), .B (n_5375), .C (n_3544), .D (n_5376), .Q
       (n_3993));
  AN22X1 g41054(.A (n_3538), .B (n_5377), .C (n_3540), .D (n_5378), .Q
       (n_3992));
  AN22X1 g41055(.A (n_3536), .B (n_5383), .C (n_3546), .D (n_5384), .Q
       (n_3991));
  AN22X1 g41056(.A (n_3547), .B (n_5385), .C (n_3504), .D (n_5386), .Q
       (n_3990));
  AN22X1 g41057(.A (n_3542), .B (n_5530), .C (n_3544), .D (n_5531), .Q
       (n_3989));
  AN22X1 g41058(.A (n_3538), .B (n_5532), .C (n_3540), .D (n_5533), .Q
       (n_3988));
  AN22X1 g41059(.A (n_3548), .B (n_4852), .C (n_3557), .D (n_4853), .Q
       (n_3987));
  AN22X1 g41060(.A (n_6768), .B (n_4854), .C (n_6767), .D (n_4855), .Q
       (n_3986));
  AN22X1 g41061(.A (n_6768), .B (n_5102), .C (n_6767), .D (n_5103), .Q
       (n_3985));
  AN22X1 g41062(.A (n_3548), .B (n_5100), .C (n_3557), .D (n_5101), .Q
       (n_3984));
  AN22X1 g41063(.A (n_3553), .B (n_5094), .C (n_3554), .D (n_5095), .Q
       (n_3983));
  AN22X1 g41064(.A (n_3549), .B (n_5092), .C (n_3551), .D (n_5093), .Q
       (n_3982));
  AN22X1 g41065(.A (n_3553), .B (n_4846), .C (n_3554), .D (n_4847), .Q
       (n_3981));
  AN22X1 g41066(.A (n_3301), .B (n_5419), .C (n_3512), .D (n_5420), .Q
       (n_3980));
  AN22X1 g41067(.A (n_3522), .B (n_4749), .C (n_3507), .D (n_4748), .Q
       (n_3979));
  AN22X1 g41068(.A (n_6768), .B (n_5536), .C (n_6767), .D (n_5537), .Q
       (n_3978));
  AN22X1 g41069(.A (n_3553), .B (n_5373), .C (n_3554), .D (n_5374), .Q
       (n_3977));
  AN22X1 g41070(.A (n_3549), .B (n_5371), .C (n_3551), .D (n_5372), .Q
       (n_3976));
  AN22X1 g41071(.A (n_6768), .B (n_5381), .C (n_6767), .D (n_5382), .Q
       (n_3975));
  AN22X1 g41072(.A (n_3548), .B (n_5379), .C (n_3557), .D (n_5380), .Q
       (n_3974));
  AN22X1 g41073(.A (n_3553), .B (n_5528), .C (n_3554), .D (n_5529), .Q
       (n_3973));
  AN22X1 g41074(.A (n_3549), .B (n_5526), .C (n_3551), .D (n_5527), .Q
       (n_3972));
  AO22X1 g41075(.A (n_3536), .B (n_5228), .C (n_3546), .D (n_5229), .Q
       (n_3971));
  AN22X1 g41077(.A (n_3542), .B (n_5158), .C (n_3544), .D (n_5159), .Q
       (n_3969));
  AO22X1 g41078(.A (n_3538), .B (n_5160), .C (n_3540), .D (n_5161), .Q
       (n_3968));
  AO22X1 g41079(.A (n_3536), .B (n_5166), .C (n_3546), .D (n_5167), .Q
       (n_3967));
  AO22X1 g41080(.A (n_3547), .B (n_5168), .C (n_3504), .D (n_5169), .Q
       (n_3966));
  AO22X1 g41081(.A (n_3536), .B (n_5073), .C (n_3546), .D (n_5074), .Q
       (n_3965));
  AO22X1 g41083(.A (n_3547), .B (n_5075), .C (n_3504), .D (n_5076), .Q
       (n_3963));
  AO22X1 g41084(.A (n_3538), .B (n_5501), .C (n_3540), .D (n_5502), .Q
       (n_3962));
  AO22X1 g41086(.A (n_3538), .B (n_5067), .C (n_3540), .D (n_5068), .Q
       (n_3960));
  AO22X1 g41088(.A (n_3547), .B (n_5509), .C (n_3504), .D (n_5510), .Q
       (n_3958));
  NO2X1 g41089(.A (n_3657), .B (n_3658), .Q (n_3957));
  AO22X1 g41090(.A (n_3538), .B (n_5005), .C (n_3540), .D (n_5006), .Q
       (n_3956));
  AN22X1 g41091(.A (n_3536), .B (n_5011), .C (n_3546), .D (n_5012), .Q
       (n_3955));
  AN22X1 g41092(.A (n_3547), .B (n_5013), .C (n_3504), .D (n_5014), .Q
       (n_3954));
  AN22X1 g41093(.A (n_3536), .B (n_4980), .C (n_3546), .D (n_4981), .Q
       (n_3953));
  AN22X1 g41094(.A (n_3547), .B (n_4982), .C (n_3504), .D (n_4983), .Q
       (n_3952));
  AN22X1 g41096(.A (n_3538), .B (n_4974), .C (n_3540), .D (n_4975), .Q
       (n_3950));
  AO22X1 g41097(.A (n_3542), .B (n_4910), .C (n_3544), .D (n_4911), .Q
       (n_3949));
  AN22X1 g41098(.A (n_3538), .B (n_4912), .C (n_3540), .D (n_4913), .Q
       (n_3948));
  AO22X1 g41100(.A (n_3547), .B (n_4920), .C (n_3504), .D (n_4921), .Q
       (n_3946));
  AN22X1 g41101(.A (n_3536), .B (n_5414), .C (n_3546), .D (n_5415), .Q
       (n_3945));
  AN22X1 g41102(.A (n_3547), .B (n_5416), .C (n_3504), .D (n_5417), .Q
       (n_3944));
  AN22X1 g41103(.A (n_3542), .B (n_5406), .C (n_3544), .D (n_5407), .Q
       (n_3943));
  AN22X1 g41104(.A (n_3538), .B (n_5408), .C (n_3540), .D (n_5409), .Q
       (n_3942));
  AN22X1 g41107(.A (n_3536), .B (n_5290), .C (n_3546), .D (n_5291), .Q
       (n_3939));
  AN22X1 g41108(.A (n_3547), .B (n_5292), .C (n_3504), .D (n_5293), .Q
       (n_3938));
  NA2X1 g41109(.A (n_3653), .B (n_3654), .Q (n_3937));
  NA2X1 g41111(.A (n_3649), .B (n_3650), .Q (n_3935));
  AO22X1 g41114(.A (n_3538), .B (n_5222), .C (n_3540), .D (n_5223), .Q
       (n_3932));
  AO22X1 g41116(.A (n_3548), .B (n_5224), .C (n_3557), .D (n_5225), .Q
       (n_3930));
  AN22X1 g41117(.A (n_3553), .B (n_5156), .C (n_3554), .D (n_5157), .Q
       (n_3929));
  NA2X1 g41123(.A (n_3634), .B (n_3633), .Q (n_3923));
  AO22X1 g41126(.A (n_3553), .B (n_5063), .C (n_3554), .D (n_5064), .Q
       (n_3920));
  AO22X1 g41127(.A (n_6768), .B (n_5505), .C (n_6767), .D (n_5506), .Q
       (n_3919));
  NO2X1 g41129(.A (n_3625), .B (n_3626), .Q (n_3917));
  AN22X1 g41131(.A (n_3548), .B (n_5007), .C (n_3557), .D (n_5008), .Q
       (n_3915));
  AN22X1 g41132(.A (n_6768), .B (n_5009), .C (n_6767), .D (n_5010), .Q
       (n_3914));
  AN22X1 g41133(.A (n_6768), .B (n_4978), .C (n_6767), .D (n_4979), .Q
       (n_3913));
  AN22X1 g41134(.A (n_3548), .B (n_4976), .C (n_3557), .D (n_4977), .Q
       (n_3912));
  NA2X1 g41135(.A (n_3622), .B (n_3621), .Q (n_3911));
  AN22X1 g41136(.A (n_3549), .B (n_4968), .C (n_3551), .D (n_4969), .Q
       (n_3910));
  NA2X1 g41137(.A (n_3620), .B (n_3619), .Q (n_3909));
  AN22X1 g41138(.A (n_3553), .B (n_4908), .C (n_3554), .D (n_4909), .Q
       (n_3908));
  NA2X1 g41139(.A (n_3618), .B (n_3617), .Q (n_3907));
  AN22X1 g41141(.A (n_6768), .B (n_5412), .C (n_6767), .D (n_5413), .Q
       (n_3905));
  AN22X1 g41142(.A (n_3548), .B (n_5410), .C (n_3557), .D (n_5411), .Q
       (n_3904));
  AN22X1 g41143(.A (n_3549), .B (n_5402), .C (n_3551), .D (n_5403), .Q
       (n_3903));
  AN22X1 g41144(.A (n_3553), .B (n_5404), .C (n_3554), .D (n_5405), .Q
       (n_3902));
  NA2X1 g41145(.A (n_3613), .B (n_3614), .Q (n_3901));
  NA2X1 g41146(.A (n_3612), .B (n_3611), .Q (n_3900));
  NA2X1 g41147(.A (n_3610), .B (n_3609), .Q (n_3899));
  NA2X1 g41149(.A (n_3607), .B (n_3608), .Q (n_3897));
  NA2X1 g41151(.A (n_3603), .B (n_3604), .Q (n_3895));
  AO22X1 g41153(.A (n_3549), .B (n_5216), .C (n_3551), .D (n_5217), .Q
       (n_3893));
  AN22X1 g41155(.A (n_3524), .B (n_4557), .C (n_3514), .D (n_4558), .Q
       (n_3891));
  AN22X1 g41156(.A (n_3516), .B (n_4551), .C (n_3512), .D (n_4552), .Q
       (n_3890));
  NA2X1 g41158(.A (n_3600), .B (n_3595), .Q (n_3888));
  AO22X1 g41160(.A (n_3296), .B (n_4564), .C (n_3509), .D (n_4556), .Q
       (n_3886));
  AN22X1 g41161(.A (n_3524), .B (n_4929), .C (n_3514), .D (n_4930), .Q
       (n_3885));
  AN22X1 g41162(.A (n_3301), .B (n_4923), .C (n_3512), .D (n_4924), .Q
       (n_3884));
  AN22X1 g41163(.A (n_3295), .B (n_4936), .C (n_3505), .D (n_4922), .Q
       (n_3883));
  AN22X1 g41164(.A (n_3510), .B (n_4927), .C (n_3526), .D (n_4926), .Q
       (n_3882));
  AO22X1 g41165(.A (n_3509), .B (n_4928), .C (n_3305), .D (n_4933), .Q
       (n_3881));
  AO22X1 g41167(.A (n_3518), .B (n_4683), .C (n_3517), .D (n_4684), .Q
       (n_3879));
  AN22X1 g41168(.A (n_3524), .B (n_4681), .C (n_3514), .D (n_4682), .Q
       (n_3878));
  AN22X1 g41169(.A (n_3301), .B (n_4675), .C (n_3512), .D (n_4676), .Q
       (n_3877));
  AO22X1 g41171(.A (n_3510), .B (n_4679), .C (n_3509), .D (n_4680), .Q
       (n_3875));
  AO22X1 g41172(.A (n_3296), .B (n_4688), .C (n_3526), .D (n_4678), .Q
       (n_3874));
  AN22X1 g41174(.A (n_3524), .B (n_4650), .C (n_3514), .D (n_4651), .Q
       (n_3872));
  AN22X1 g41175(.A (n_3301), .B (n_4644), .C (n_3512), .D (n_4645), .Q
       (n_3871));
  AO22X1 g41177(.A (n_3296), .B (n_4657), .C (n_3526), .D (n_4647), .Q
       (n_3869));
  AO22X1 g41178(.A (n_3510), .B (n_4648), .C (n_3509), .D (n_4649), .Q
       (n_3868));
  NA2X1 g41180(.A (n_3579), .B (n_3580), .Q (n_3866));
  AO22X1 g41183(.A (n_3547), .B (n_4579), .C (n_3504), .D (n_4580), .Q
       (n_3863));
  AN22X1 g41184(.A (n_3542), .B (n_4941), .C (n_3544), .D (n_4942), .Q
       (n_3862));
  AN22X1 g41185(.A (n_3538), .B (n_4943), .C (n_3540), .D (n_4944), .Q
       (n_3861));
  AN22X1 g41186(.A (n_3536), .B (n_4949), .C (n_3546), .D (n_4950), .Q
       (n_3860));
  AN22X1 g41187(.A (n_3547), .B (n_4951), .C (n_3504), .D (n_4952), .Q
       (n_3859));
  AO22X1 g41188(.A (n_3542), .B (n_4693), .C (n_3544), .D (n_4694), .Q
       (n_3858));
  AN22X1 g41191(.A (n_3547), .B (n_4703), .C (n_3504), .D (n_4704), .Q
       (n_3855));
  AN22X1 g41192(.A (n_3542), .B (n_4662), .C (n_3544), .D (n_4663), .Q
       (n_3854));
  AN22X1 g41193(.A (n_3538), .B (n_4664), .C (n_3540), .D (n_4665), .Q
       (n_3853));
  AN22X1 g41194(.A (n_3536), .B (n_4670), .C (n_3546), .D (n_4671), .Q
       (n_3852));
  AN22X1 g41195(.A (n_3547), .B (n_4672), .C (n_3504), .D (n_4673), .Q
       (n_3851));
  NA2X1 g41196(.A (n_3583), .B (n_3588), .Q (n_3850));
  AN22X1 g41199(.A (n_3553), .B (n_4939), .C (n_3554), .D (n_4940), .Q
       (n_3847));
  AO22X1 g41201(.A (n_3553), .B (n_4691), .C (n_3554), .D (n_4692), .Q
       (n_3845));
  AN22X1 g41202(.A (n_3549), .B (n_4658), .C (n_3551), .D (n_4659), .Q
       (n_3844));
  AN22X1 g41203(.A (n_3553), .B (n_4660), .C (n_3554), .D (n_4661), .Q
       (n_3843));
  NA2X1 g41205(.A (n_3586), .B (n_3587), .Q (n_3841));
  AN22X1 g41206(.A (n_3548), .B (n_4945), .C (n_3557), .D (n_4946), .Q
       (n_3840));
  AN22X1 g41207(.A (n_6768), .B (n_4947), .C (n_6767), .D (n_4948), .Q
       (n_3839));
  AO22X1 g41208(.A (n_3548), .B (n_4697), .C (n_3557), .D (n_4698), .Q
       (n_3838));
  AN22X1 g41209(.A (n_6768), .B (n_4699), .C (n_6767), .D (n_4700), .Q
       (n_3837));
  AO22X1 g41210(.A (n_3548), .B (n_4666), .C (n_3557), .D (n_4667), .Q
       (n_3836));
  AN22X1 g41212(.A (n_3536), .B (n_5042), .C (n_3546), .D (n_5043), .Q
       (n_3834));
  AN22X1 g41214(.A (n_3542), .B (n_5034), .C (n_3544), .D (n_5035), .Q
       (n_3832));
  AN22X1 g41215(.A (n_3538), .B (n_5036), .C (n_3540), .D (n_5037), .Q
       (n_3831));
  AN22X1 g41216(.A (n_3542), .B (n_4817), .C (n_3544), .D (n_4818), .Q
       (n_3830));
  AN22X1 g41217(.A (n_3538), .B (n_4819), .C (n_3540), .D (n_4820), .Q
       (n_3829));
  AN22X1 g41218(.A (n_3536), .B (n_4825), .C (n_3546), .D (n_4826), .Q
       (n_3828));
  AN22X1 g41219(.A (n_3547), .B (n_4827), .C (n_3504), .D (n_4828), .Q
       (n_3827));
  AN22X1 g41220(.A (n_6768), .B (n_5040), .C (n_6767), .D (n_5041), .Q
       (n_3826));
  AO22X1 g41221(.A (n_3548), .B (n_5038), .C (n_3557), .D (n_5039), .Q
       (n_3825));
  AN22X1 g41222(.A (n_3549), .B (n_5030), .C (n_3551), .D (n_5031), .Q
       (n_3824));
  AN22X1 g41223(.A (n_3553), .B (n_5032), .C (n_3554), .D (n_5033), .Q
       (n_3823));
  AN22X1 g41224(.A (n_3549), .B (n_4813), .C (n_3551), .D (n_4814), .Q
       (n_3822));
  AN22X1 g41225(.A (n_3553), .B (n_4815), .C (n_3554), .D (n_4816), .Q
       (n_3821));
  AN22X1 g41226(.A (n_3548), .B (n_4821), .C (n_3557), .D (n_4822), .Q
       (n_3820));
  AN22X1 g41227(.A (n_6768), .B (n_4823), .C (n_6767), .D (n_4824), .Q
       (n_3819));
  AN22X1 g41228(.A (n_3301), .B (n_5016), .C (n_3512), .D (n_5017), .Q
       (n_3818));
  AN22X1 g41229(.A (n_3296), .B (n_5029), .C (n_3505), .D (n_5015), .Q
       (n_3817));
  AN22X1 g41230(.A (n_3510), .B (n_5020), .C (n_3526), .D (n_5019), .Q
       (n_3816));
  AN22X1 g41231(.A (n_3301), .B (n_4799), .C (n_3512), .D (n_4800), .Q
       (n_3815));
  AN22X1 g41232(.A (n_3296), .B (n_4812), .C (n_3505), .D (n_4798), .Q
       (n_3814));
  AN22X1 g41233(.A (n_3510), .B (n_4803), .C (n_3526), .D (n_4802), .Q
       (n_3813));
  AN22X1 g41234(.A (n_3524), .B (n_5022), .C (n_3514), .D (n_5023), .Q
       (n_3812));
  AN22X1 g41235(.A (n_3509), .B (n_5021), .C (n_3305), .D (n_5026), .Q
       (n_3811));
  AN22X1 g41236(.A (n_3522), .B (n_5028), .C (n_3298), .D (n_5027), .Q
       (n_3810));
  AO22X2 g41237(.A (n_3518), .B (n_4807), .C (n_3517), .D (n_4808), .Q
       (n_3809));
  AN22X1 g41238(.A (n_3524), .B (n_4805), .C (n_3514), .D (n_4806), .Q
       (n_3808));
  AN22X1 g41239(.A (n_3509), .B (n_4804), .C (n_3305), .D (n_4809), .Q
       (n_3807));
  AN22X1 g41240(.A (n_3522), .B (n_4811), .C (n_3298), .D (n_4810), .Q
       (n_3806));
  ON22X1 g41244(.A (n_3537), .B (n_3360), .C (n_3539), .D (n_3368), .Q
       (n_3802));
  AN22X1 g41245(.A (n_6768), .B (n_4885), .C (n_6767), .D (n_4886), .Q
       (n_3801));
  AN22X1 g41246(.A (n_3548), .B (n_4883), .C (n_3557), .D (n_4884), .Q
       (n_3800));
  AO22X2 g41247(.A (n_3553), .B (n_4753), .C (n_3554), .D (n_4754), .Q
       (n_3799));
  AN22X1 g41248(.A (n_3548), .B (n_4790), .C (n_3557), .D (n_4791), .Q
       (n_3798));
  AN22X1 g41249(.A (n_6768), .B (n_4792), .C (n_6767), .D (n_4793), .Q
       (n_3797));
  AN22X1 g41250(.A (n_3549), .B (n_4782), .C (n_3551), .D (n_4783), .Q
       (n_3796));
  AN22X1 g41251(.A (n_3542), .B (n_4786), .C (n_3544), .D (n_4787), .Q
       (n_3795));
  AN22X1 g41252(.A (n_3538), .B (n_4788), .C (n_3540), .D (n_4789), .Q
       (n_3794));
  AN22X1 g41253(.A (n_3548), .B (n_4759), .C (n_3557), .D (n_4760), .Q
       (n_3793));
  AN22X1 g41254(.A (n_6768), .B (n_4761), .C (n_6767), .D (n_4762), .Q
       (n_3792));
  NA2X1 g41255(.A (n_3570), .B (n_3569), .Q (n_3791));
  NA2X1 g41256(.A (n_3574), .B (n_3575), .Q (n_3790));
  AO22X1 g41257(.A (n_3538), .B (n_4757), .C (n_3540), .D (n_4758), .Q
       (n_3789));
  AN22X1 g41258(.A (n_3553), .B (n_4784), .C (n_3554), .D (n_4785), .Q
       (n_3788));
  AN22X1 g41259(.A (n_3536), .B (n_4887), .C (n_3546), .D (n_4888), .Q
       (n_3787));
  AN22X1 g41260(.A (n_3547), .B (n_4889), .C (n_3504), .D (n_4890), .Q
       (n_3786));
  AO22X2 g41262(.A (n_3547), .B (n_4796), .C (n_3504), .D (n_4797), .Q
       (n_3784));
  NO2X1 g41263(.A (n_3566), .B (n_3565), .Q (n_3783));
  AN22X1 g41264(.A (n_3547), .B (n_4765), .C (n_3504), .D (n_4766), .Q
       (n_3782));
  AN22X1 g41265(.A (n_3516), .B (n_4861), .C (n_3512), .D (n_4862), .Q
       (n_3781));
  AN22X1 g41266(.A (n_3510), .B (n_4865), .C (n_3526), .D (n_4864), .Q
       (n_3780));
  AN22X1 g41267(.A (n_3509), .B (n_4866), .C (n_3303), .D (n_4871), .Q
       (n_3779));
  AN22X1 g41268(.A (n_3516), .B (n_4737), .C (n_3512), .D (n_4738), .Q
       (n_3778));
  AN22X1 g41269(.A (n_3516), .B (n_4768), .C (n_3512), .D (n_4769), .Q
       (n_3777));
  AN22X1 g41270(.A (n_3510), .B (n_4772), .C (n_3526), .D (n_4771), .Q
       (n_3776));
  AN22X1 g41271(.A (n_3509), .B (n_4773), .C (n_3303), .D (n_4778), .Q
       (n_3775));
  AN22X1 g41272(.A (n_3510), .B (n_4741), .C (n_3526), .D (n_4740), .Q
       (n_3774));
  AN22X1 g41273(.A (n_3509), .B (n_4742), .C (n_3303), .D (n_4747), .Q
       (n_3773));
  AN22X1 g41274(.A (n_3524), .B (n_4867), .C (n_3514), .D (n_4868), .Q
       (n_3772));
  AN22X1 g41275(.A (n_3296), .B (n_4874), .C (n_3505), .D (n_4860), .Q
       (n_3771));
  AN22X1 g41276(.A (n_3522), .B (n_4873), .C (n_3507), .D (n_4872), .Q
       (n_3770));
  ON22X1 g41277(.A (n_3519), .B (n_3367), .C (n_3302), .D (n_3378), .Q
       (n_3769));
  AN22X1 g41278(.A (n_3524), .B (n_4774), .C (n_3514), .D (n_4775), .Q
       (n_3768));
  AN22X1 g41279(.A (n_3296), .B (n_4781), .C (n_3505), .D (n_4767), .Q
       (n_3767));
  AN22X1 g41280(.A (n_3522), .B (n_4780), .C (n_3507), .D (n_4779), .Q
       (n_3766));
  AN22X1 g41281(.A (n_3524), .B (n_4743), .C (n_3514), .D (n_4744), .Q
       (n_3765));
  AN22X1 g41282(.A (n_3296), .B (n_4750), .C (n_3505), .D (n_4736), .Q
       (n_3764));
  AN22X1 g41283(.A (n_3548), .B (n_5534), .C (n_3557), .D (n_5535), .Q
       (n_3763));
  NA2X1 g41284(.A (n_3512), .B (n_5327), .Q (n_3762));
  NA2X1 g41285(.A (n_3301), .B (n_5326), .Q (n_3761));
  NO2I1X1 g41288(.B (n_3302), .AN (n_5335), .Q (n_3758));
  NO2I1X1 g41291(.B (n_3302), .AN (n_5304), .Q (n_3755));
  NO2I1X1 g41292(.B (n_3302), .AN (n_4591), .Q (n_3754));
  NA2X1 g41293(.A (n_3301), .B (n_4706), .Q (n_3753));
  NA2X1 g41294(.A (n_3512), .B (n_4707), .Q (n_3752));
  NO2I1X1 g41295(.B (n_3506), .AN (n_4705), .Q (n_3751));
  NO2I1X1 g41296(.B (n_3302), .AN (n_4715), .Q (n_3750));
  NO2I1X1 g41297(.B (n_3519), .AN (n_4714), .Q (n_3749));
  NO2I1X1 g41299(.B (n_3302), .AN (n_5459), .Q (n_3747));
  NO2I1X1 g41301(.B (n_3302), .AN (n_4622), .Q (n_3745));
  NO2I1X1 g41302(.B (n_3297), .AN (n_4717), .Q (n_3744));
  NA2X1 g41303(.A (n_3505), .B (n_4829), .Q (n_3743));
  NA2X1 g41307(.A (n_3526), .B (n_4833), .Q (n_3739));
  NA2X1 g41308(.A (n_3510), .B (n_4834), .Q (n_3738));
  NA2X1 g41309(.A (n_3505), .B (n_5511), .Q (n_3737));
  NO2I1X1 g41310(.B (n_3302), .AN (n_4839), .Q (n_3736));
  NO2I1X1 g41311(.B (n_3519), .AN (n_4838), .Q (n_3735));
  NA2X1 g41312(.A (n_3524), .B (n_4836), .Q (n_3734));
  NA2X1 g41313(.A (n_3514), .B (n_4837), .Q (n_3733));
  NO2I1X1 g41318(.B (n_3302), .AN (n_5521), .Q (n_3728));
  NO2I1X1 g41319(.B (n_3519), .AN (n_5520), .Q (n_3727));
  NO2I1X1 g41322(.B (n_3302), .AN (n_5366), .Q (n_3724));
  NA2X1 g41325(.A (n_3296), .B (n_4843), .Q (n_3721));
  NA2X1 g41327(.A (n_3296), .B (n_5525), .Q (n_3719));
  NA2X1 g41330(.A (n_3517), .B (n_5149), .Q (n_3716));
  NA2X1 g41331(.A (n_3518), .B (n_5148), .Q (n_3715));
  NO2I1X1 g41332(.B (n_3515), .AN (n_5147), .Q (n_3714));
  NO2I1X1 g41333(.B (n_3525), .AN (n_5146), .Q (n_3713));
  NO2I1X1 g41334(.B (n_3513), .AN (n_5141), .Q (n_3712));
  NO2I1X1 g41335(.B (n_3300), .AN (n_5140), .Q (n_3711));
  NO2I1X1 g41336(.B (n_3506), .AN (n_5139), .Q (n_3710));
  NO2I1X1 g41337(.B (n_3302), .AN (n_4994), .Q (n_3709));
  NO2I1X1 g41338(.B (n_3519), .AN (n_4993), .Q (n_3708));
  NA2X1 g41339(.A (n_3514), .B (n_4961), .Q (n_3707));
  NA2X1 g41340(.A (n_3524), .B (n_4960), .Q (n_3706));
  NO2I1X1 g41341(.B (n_3525), .AN (n_4898), .Q (n_3705));
  NO2I1X1 g41342(.B (n_3515), .AN (n_4899), .Q (n_3704));
  NO2I1X1 g41343(.B (n_3302), .AN (n_5273), .Q (n_3703));
  NO2I1X1 g41344(.B (n_3506), .AN (n_5263), .Q (n_3702));
  NA2X1 g41345(.A (n_3517), .B (n_5242), .Q (n_3701));
  NA2X1 g41346(.A (n_3518), .B (n_5241), .Q (n_3700));
  NO2I1X1 g41347(.B (n_3515), .AN (n_5240), .Q (n_3699));
  NO2I1X1 g41348(.B (n_3525), .AN (n_5239), .Q (n_3698));
  NO2I1X1 g41349(.B (n_3513), .AN (n_5234), .Q (n_3697));
  NO2I1X1 g41350(.B (n_3300), .AN (n_5233), .Q (n_3696));
  NO2I1X1 g41351(.B (n_3506), .AN (n_5232), .Q (n_3695));
  NO2I1X1 g41352(.B (n_3302), .AN (n_5211), .Q (n_3694));
  NO2I1X1 g41353(.B (n_3519), .AN (n_5210), .Q (n_3693));
  NA2X1 g41354(.A (n_3520), .B (n_5142), .Q (n_3692));
  NO2I1X1 g41355(.B (n_3294), .AN (n_5153), .Q (n_3691));
  NO2I1X1 g41356(.B (n_3527), .AN (n_5143), .Q (n_3690));
  NO2I1X1 g41357(.B (n_3511), .AN (n_5144), .Q (n_3689));
  NO2I1X1 g41359(.B (n_3299), .AN (n_5145), .Q (n_3688));
  NO2I1X1 g41360(.B (n_3297), .AN (n_5151), .Q (n_3687));
  NO2I1X1 g41361(.B (n_3523), .AN (n_5152), .Q (n_3686));
  NO2I1X1 g41364(.B (n_3294), .AN (n_5060), .Q (n_3683));
  NA2X1 g41365(.A (n_3305), .B (n_5491), .Q (n_3682));
  NA2X1 g41366(.A (n_3509), .B (n_5486), .Q (n_3681));
  NO2I1X1 g41369(.B (n_3521), .AN (n_4956), .Q (n_3678));
  NO2I1X1 g41370(.B (n_3294), .AN (n_5277), .Q (n_3677));
  NO2I1X1 g41371(.B (n_3527), .AN (n_5267), .Q (n_3676));
  NO2I1X1 g41372(.B (n_3511), .AN (n_5268), .Q (n_3675));
  NO2I1X1 g41373(.B (n_3304), .AN (n_5274), .Q (n_3674));
  NO2I1X1 g41374(.B (n_3299), .AN (n_5269), .Q (n_3673));
  NO2I1X1 g41375(.B (n_3297), .AN (n_5275), .Q (n_3672));
  NO2I1X1 g41376(.B (n_3523), .AN (n_5276), .Q (n_3671));
  NA2X1 g41377(.A (n_3520), .B (n_5235), .Q (n_3670));
  NO2I1X1 g41378(.B (n_3294), .AN (n_5246), .Q (n_3669));
  NO2I1X1 g41379(.B (n_3297), .AN (n_5244), .Q (n_3668));
  NO2I1X1 g41380(.B (n_3523), .AN (n_5245), .Q (n_3667));
  NO2I1X1 g41381(.B (n_3527), .AN (n_5236), .Q (n_3666));
  NO2I1X1 g41382(.B (n_3511), .AN (n_5237), .Q (n_3665));
  NO2I1X1 g41383(.B (n_3304), .AN (n_5243), .Q (n_3664));
  NO2I1X1 g41384(.B (n_3299), .AN (n_5238), .Q (n_3663));
  NO2I1X1 g41389(.B (n_3543), .AN (n_5004), .Q (n_3658));
  NO2I1X1 g41390(.B (n_3541), .AN (n_5003), .Q (n_3657));
  NA2X1 g41393(.A (n_3544), .B (n_5252), .Q (n_3654));
  NA2X1 g41394(.A (n_3542), .B (n_5251), .Q (n_3653));
  NA2X1 g41397(.A (n_3546), .B (n_5260), .Q (n_3650));
  NA2X1 g41398(.A (n_3536), .B (n_5259), .Q (n_3649));
  NA2X1 g41413(.A (n_3554), .B (n_5498), .Q (n_3634));
  NA2X1 g41414(.A (n_3553), .B (n_5497), .Q (n_3633));
  NO2I1X1 g41421(.B (n_3552), .AN (n_5000), .Q (n_3626));
  NO2I1X1 g41422(.B (n_3550), .AN (n_4999), .Q (n_3625));
  NA2X1 g41425(.A (n_3554), .B (n_4971), .Q (n_3622));
  NA2X1 g41426(.A (n_3553), .B (n_4970), .Q (n_3621));
  NA2X1 g41427(.A (n_3551), .B (n_4907), .Q (n_3620));
  NA2X1 g41428(.A (n_3549), .B (n_4906), .Q (n_3619));
  NA2X1 g41429(.A (n_6767), .B (n_4917), .Q (n_3618));
  NA2X1 g41430(.A (n_6768), .B (n_4916), .Q (n_3617));
  NA2X1 g41433(.A (n_3551), .B (n_5279), .Q (n_3614));
  NA2X1 g41434(.A (n_3549), .B (n_5278), .Q (n_3613));
  NA2X1 g41435(.A (n_3554), .B (n_5281), .Q (n_3612));
  NA2X1 g41436(.A (n_3553), .B (n_5280), .Q (n_3611));
  NA2X1 g41437(.A (n_3557), .B (n_5287), .Q (n_3610));
  NA2X1 g41438(.A (n_3548), .B (n_5286), .Q (n_3609));
  NA2X1 g41439(.A (n_3551), .B (n_5248), .Q (n_3608));
  NA2X1 g41440(.A (n_3549), .B (n_5247), .Q (n_3607));
  NA2X1 g41443(.A (n_3557), .B (n_5256), .Q (n_3604));
  NA2X1 g41444(.A (n_3548), .B (n_5255), .Q (n_3603));
  NA2X1 g41448(.A (n_3510), .B (n_4555), .Q (n_3600));
  NO2X1 g41449(.A (n_3521), .B (n_3366), .Q (n_3599));
  NA2X1 g41454(.A (n_3507), .B (n_4562), .Q (n_3595));
  AND2X1 g41457(.A (n_3517), .B (n_4653), .Q (n_3592));
  NO2I1X1 g41460(.B (n_3521), .AN (n_4801), .Q (n_3589));
  NA2X1 g41461(.A (n_3551), .B (n_4566), .Q (n_3588));
  NA2X1 g41462(.A (n_6767), .B (n_4576), .Q (n_3587));
  NA2X1 g41463(.A (n_6768), .B (n_4575), .Q (n_3586));
  NA2X1 g41466(.A (n_3549), .B (n_4565), .Q (n_3583));
  NA2X1 g41469(.A (n_3544), .B (n_4570), .Q (n_3580));
  NA2X1 g41470(.A (n_3542), .B (n_4569), .Q (n_3579));
  NA2X1 g41474(.A (n_3551), .B (n_4752), .Q (n_3575));
  NA2X1 g41475(.A (n_3549), .B (n_4751), .Q (n_3574));
  NA2X1 g41479(.A (n_3542), .B (n_4755), .Q (n_3570));
  NA2X1 g41480(.A (n_3544), .B (n_4756), .Q (n_3569));
  NO2I1X1 g41483(.B (n_3535), .AN (n_4763), .Q (n_3566));
  NO2I1X1 g41484(.B (n_3545), .AN (n_4764), .Q (n_3565));
  NO2I1X1 g41485(.B (n_3521), .AN (n_4739), .Q (n_3564));
  NO2I1X1 g41486(.B (n_3521), .AN (n_4770), .Q (n_3563));
  NO2I1X1 g41487(.B (n_3521), .AN (n_4863), .Q (n_3562));
  AND2X2 g41488(.A (n_3517), .B (n_4870), .Q (n_3561));
  NO2I1X1 g41489(.B (n_3519), .AN (n_4869), .Q (n_3560));
  NO2I1X1 g41490(.B (n_3519), .AN (n_4745), .Q (n_3559));
  NO2I1X1 g41491(.B (n_3302), .AN (n_4746), .Q (n_3558));
  INX4 g41492(.A (n_3534), .Q (n_3557));
  INX4 g41495(.A (n_3531), .Q (n_3554));
  INX6 g41496(.A (n_3530), .Q (n_3553));
  INX4 g41497(.A (n_3552), .Q (n_3551));
  INX8 g41498(.A (n_3550), .Q (n_3549));
  INX6 g41499(.A (n_3529), .Q (n_3548));
  INX8 g41500(.A (n_3528), .Q (n_3547));
  INX4 g41501(.A (n_3545), .Q (n_3546));
  INX8 g41502(.A (n_3543), .Q (n_3544));
  INX8 g41503(.A (n_3541), .Q (n_3542));
  INX4 g41504(.A (n_3539), .Q (n_3540));
  INX6 g41505(.A (n_3537), .Q (n_3538));
  INX4 g41506(.A (n_3535), .Q (n_3536));
  NA2X2 g41507(.A (n_3500), .B (n_3485), .Q (n_3534));
  NA2X4 g41510(.A (n_3500), .B (n_3482), .Q (n_3531));
  NA2X4 g41511(.A (n_3500), .B (n_3293), .Q (n_3530));
  NA2X4 g41512(.A (n_3500), .B (n_3292), .Q (n_3552));
  NA2X4 g41513(.A (n_3500), .B (n_3491), .Q (n_3550));
  NA2X2 g41514(.A (n_3500), .B (n_3484), .Q (n_3529));
  NA2X4 g41515(.A (n_3498), .B (n_3291), .Q (n_3528));
  NA2X2 g41516(.A (n_3498), .B (n_3485), .Q (n_3545));
  NA2X4 g41517(.A (n_3498), .B (n_3292), .Q (n_3543));
  NA2X4 g41518(.A (n_3498), .B (n_3491), .Q (n_3541));
  NA2X4 g41519(.A (n_3498), .B (n_3482), .Q (n_3539));
  NA2X4 g41520(.A (n_3498), .B (n_3293), .Q (n_3537));
  NA2X2 g41521(.A (n_3498), .B (n_3484), .Q (n_3535));
  INX4 g41531(.A (n_3527), .Q (n_3526));
  INX4 g41532(.A (n_3525), .Q (n_3524));
  INX8 g41533(.A (n_3523), .Q (n_3522));
  INX4 g41534(.A (n_3521), .Q (n_3520));
  INX6 g41535(.A (n_3519), .Q (n_3518));
  INX4 g41549(.A (n_3515), .Q (n_3514));
  INX4 g41550(.A (n_3513), .Q (n_3512));
  INX6 g41551(.A (n_3511), .Q (n_3510));
  INX1 g41554(.A (n_3299), .Q (n_3508));
  INX1 g41556(.A (n_3509), .Q (n_3299));
  INX2 g41575(.A (n_3294), .Q (n_3295));
  INX6 g41580(.A (n_3506), .Q (n_3505));
  INX6 g41581(.A (n_3503), .Q (n_3504));
  AND2X4 g41582(.A (n_3499), .B (n_3484), .Q (n_3305));
  OR2X4 g41584(.A (n_3282), .B (n_3488), .Q (n_3527));
  OR2X4 g41585(.A (n_3502), .B (n_3483), .Q (n_3525));
  OR2X4 g41586(.A (n_3282), .B (n_3486), .Q (n_3523));
  OR2X4 g41587(.A (n_3282), .B (n_3490), .Q (n_3521));
  OR2X4 g41588(.A (n_3502), .B (n_3486), .Q (n_3519));
  NA2X4 g41589(.A (n_3501), .B (n_3487), .Q (n_3302));
  AND2X4 g41590(.A (n_3501), .B (n_3487), .Q (n_3517));
  AND2X4 g41591(.A (n_3501), .B (n_3293), .Q (n_3301));
  OR2X4 g41593(.A (n_3502), .B (n_3478), .Q (n_3515));
  OR2X4 g41594(.A (n_3502), .B (n_3481), .Q (n_3513));
  OR2X4 g41595(.A (n_3282), .B (n_3489), .Q (n_3511));
  AND2X4 g41596(.A (n_3499), .B (n_3482), .Q (n_3509));
  AND2X4 g41597(.A (n_3499), .B (n_3485), .Q (n_3298));
  AND2X2 g41598(.A (n_3499), .B (n_3485), .Q (n_3507));
  AND2X4 g41599(.A (n_3499), .B (n_3487), .Q (n_3296));
  OR2X4 g41600(.A (n_3502), .B (n_3488), .Q (n_3506));
  NA2X4 g41601(.A (n_3498), .B (n_3487), .Q (n_3503));
  AO21X1 g41603(.A (n_6623), .B (instruction[22]), .C (n_3471), .Q
       (n_6011));
  AO21X1 g41605(.A (n_6623), .B (instruction[23]), .C (n_3472), .Q
       (n_6010));
  INX2 g41606(.A (n_3502), .Q (n_3501));
  INX3 g41607(.A (n_3282), .Q (n_3499));
  OR2X4 g41608(.A (n_3495), .B (n_3454), .Q (n_3502));
  AND2X4 g41609(.A (n_3495), .B (n_3458), .Q (n_3500));
  AND2X4 g41611(.A (n_3495), .B (n_3454), .Q (n_3498));
  AO21X1 g41614(.A (n_3480), .B (instruction[16]), .C (n_3493), .Q
       (n_6004));
  AO21X1 g41615(.A (n_3480), .B (instruction[18]), .C (n_3493), .Q
       (n_6002));
  AO221X1 g41616(.A (\instruction[7]_39562 ), .B (branch_type), .C
       (jal_type), .D (n_6723), .E (n_3496), .Q (n_6013));
  AO21X1 g41617(.A (n_3480), .B (instruction[15]), .C (n_3493), .Q
       (n_6005));
  AO21X1 g41618(.A (n_3480), .B (\instruction[14]_40077 ), .C (n_3493),
       .Q (n_6006));
  AO21X1 g41619(.A (n_3480), .B (instruction[19]), .C (n_3493), .Q
       (n_6001));
  AO21X1 g41620(.A (n_3480), .B (n_6720), .C (n_3493), .Q (n_6008));
  AO21X1 g41621(.A (n_3480), .B (n_6721), .C (n_3493), .Q (n_6007));
  AO21X1 g41622(.A (n_3480), .B (instruction[17]), .C (n_3493), .Q
       (n_6003));
  NA2X2 g41623(.A (n_3281), .B (n_3473), .Q (n_6014));
  NO2X1 g41624(.A (n_3492), .B (branch_type), .Q (n_3496));
  NO2I1X4 g41627(.B (n_3479), .AN (n_6606), .Q (n_3495));
  INX1 g41629(.A (n_3493), .Q (n_3492));
  AO21X1 g41630(.A (n_3456), .B (instruction[23]), .C (n_3475), .Q
       (n_6000));
  AO21X1 g41631(.A (n_3456), .B (instruction[29]), .C (n_3475), .Q
       (n_5994));
  AO21X1 g41632(.A (n_3456), .B (instruction[24]), .C (n_3475), .Q
       (n_5999));
  AO21X1 g41633(.A (n_3456), .B (instruction[28]), .C (n_3475), .Q
       (n_5995));
  AO21X1 g41634(.A (n_3456), .B (instruction[27]), .C (n_3475), .Q
       (n_5996));
  AO21X1 g41635(.A (n_3456), .B (instruction[25]), .C (n_3475), .Q
       (n_5998));
  AO21X1 g41636(.A (n_3456), .B (n_6722), .C (n_3475), .Q (n_5993));
  AO21X1 g41637(.A (n_3456), .B (instruction[26]), .C (n_3475), .Q
       (n_5997));
  AO21X1 g41638(.A (n_3456), .B (instruction[21]), .C (n_3475), .Q
       (n_6015));
  AO21X1 g41639(.A (n_3456), .B (instruction[22]), .C (n_3475), .Q
       (n_5991));
  NA2X1 g41640(.A (n_3476), .B (n_3468), .Q (n_3494));
  NO2X1 g41641(.A (n_3474), .B (jal_type), .Q (n_3493));
  INX1 g41643(.A (n_3490), .Q (n_3491));
  INX1 g41647(.A (n_3291), .Q (n_3486));
  INX2 g41649(.A (n_3481), .Q (n_3482));
  AO21X1 g41650(.A (n_3456), .B (n_6723), .C (n_3475), .Q (n_5992));
  NO2X2 g41651(.A (n_3461), .B (n_3434), .Q (n_3479));
  NA3X2 g41652(.A (n_3446), .B (n_3434), .C (n_3435), .Q (n_6606));
  NA2X2 g41653(.A (n_3465), .B (n_3438), .Q (n_3490));
  NA2X2 g41654(.A (n_3465), .B (n_3452), .Q (n_3489));
  NA2X2 g41655(.A (n_3465), .B (n_3442), .Q (n_3488));
  AND2X4 g41656(.A (n_3477), .B (n_3455), .Q (n_3487));
  NO2X4 g41657(.A (n_3465), .B (n_3453), .Q (n_3291));
  NO2X1 g41658(.A (n_3465), .B (n_3443), .Q (n_3485));
  NA2X1 g41659(.A (n_3477), .B (n_3442), .Q (n_3478));
  OR2X2 g41660(.A (n_3465), .B (n_3439), .Q (n_3483));
  NA2X2 g41661(.A (n_3465), .B (n_3455), .Q (n_3481));
  NO2I1X1 g41662(.B (n_3476), .AN (n_3468), .Q (n_3480));
  INX1 g41663(.A (n_3465), .Q (n_3477));
  INX1 g41664(.A (n_3474), .Q (n_3475));
  AND2X1 g41665(.A (n_3467), .B (instruction[29]), .Q (n_6558));
  AND2X1 g41666(.A (n_3467), .B (n_6722), .Q (n_6559));
  AND2X1 g41667(.A (n_3467), .B (instruction[27]), .Q (n_6556));
  AND2X1 g41668(.A (n_3467), .B (instruction[28]), .Q (n_6557));
  NO2X1 g41669(.A (n_3466), .B (jal_type), .Q (n_3476));
  NA2X1 g41670(.A (n_3467), .B (n_6719), .Q (n_3474));
  AN22X1 g41671(.A (n_3290), .B (instruction[15]), .C (store_type), .D
       (\instruction[7]_39562 ), .Q (n_3473));
  AND2X1 g41672(.A (n_3467), .B (instruction[25]), .Q (n_6554));
  AO22X1 g41673(.A (n_3464), .B (\instruction[10]_39951 ), .C (n_3290),
       .D (instruction[18]), .Q (n_3472));
  AO22X1 g41674(.A (n_3464), .B (\instruction[9]_39983 ), .C (n_6453),
       .D (instruction[17]), .Q (n_3471));
  AND2X1 g41677(.A (n_3467), .B (instruction[26]), .Q (n_6555));
  NO2X1 g41679(.A (n_3464), .B (n_3290), .Q (n_3468));
  INX1 g41680(.A (n_3466), .Q (n_3467));
  NA2X1 g41681(.A (n_3462), .B (n_6561), .Q (n_3466));
  NA2I1X4 g41682(.B (n_3460), .AN (n_3459), .Q (n_3465));
  BUX6 g41687(.A (n_3290), .Q (n_6453));
  INX2 g41689(.A (n_3462), .Q (n_3290));
  OR2X2 g41690(.A (store_type), .B (branch_type), .Q (n_3464));
  NA2I1X2 g41691(.B (system_type), .AN (n_5605), .Q (n_3462));
  INX2 g41692(.A (n_3460), .Q (n_3461));
  NO2X2 g41693(.A (n_3446), .B (n_3435), .Q (n_3459));
  NA2X2 g41694(.A (n_3446), .B (n_3435), .Q (n_3460));
  INX1 g41695(.A (n_3454), .Q (n_3458));
  NO2X2 g41696(.A (n_6603), .B (n_3450), .Q (system_type));
  NO2X2 g41697(.A (n_6603), .B (n_6604), .Q (branch_type));
  INX1 g41699(.A (n_6561), .Q (n_3456));
  NO2X2 g41700(.A (n_6598), .B (n_3451), .Q (store_type));
  NO2X2 g41701(.A (n_6602), .B (n_6604), .Q (jal_type));
  NA3X2 g41702(.A (n_3449), .B (n_3447), .C (n_3444), .Q (n_6561));
  NA2X1 g41704(.A (n_3449), .B (n_3444), .Q (n_6601));
  NA3X1 g41705(.A (n_3449), .B (instruction[3]), .C (instruction[2]),
       .Q (n_6602));
  NO2X1 g41706(.A (n_3448), .B (n_3428), .Q (n_3455));
  NA2X2 g41707(.A (n_3449), .B (n_3440), .Q (n_6603));
  NO2X4 g41708(.A (n_3446), .B (n_3445), .Q (n_3454));
  INX1 g41709(.A (n_3452), .Q (n_3453));
  NA3X1 g41710(.A (instruction[4]), .B (\instruction[5]_40139 ), .C
       (n_3430), .Q (n_6599));
  NA3X1 g41711(.A (n_3431), .B (n_3437), .C (n_3430), .Q (n_3451));
  NA3X1 g41713(.A (instruction[4]), .B (instruction[6]), .C (n_3431),
       .Q (n_3450));
  NO2X2 g41714(.A (n_3448), .B (instruction[15]), .Q (n_3452));
  NA3X2 g41715(.A (instruction[6]), .B (n_3431), .C (n_3437), .Q
       (n_6604));
  NO2X2 g41716(.A (n_3441), .B (\instruction[14]_40077 ), .Q (n_6459));
  AND2X2 g41718(.A (n_6718), .B (instruction[0]), .Q (n_3449));
  NO2X1 g41719(.A (n_3438), .B (n_3433), .Q (n_3445));
  NA2X1 g41720(.A (n_3443), .B (n_3439), .Q (n_3448));
  NO2X1 g41721(.A (instruction[6]), .B (n_3437), .Q (n_3447));
  NO2X4 g41722(.A (n_3439), .B (instruction[17]), .Q (n_3446));
  INX1 g41723(.A (n_3443), .Q (n_3442));
  INX1 g41724(.A (n_5605), .Q (n_3441));
  NO2X1 g41725(.A (instruction[3]), .B (n_3436), .Q (n_3444));
  NO2X1 g41726(.A (instruction[2]), .B (instruction[3]), .Q (n_3440));
  NA2X2 g41727(.A (instruction[16]), .B (instruction[15]), .Q (n_3443));
  NO2X2 g41728(.A (n_6720), .B (n_6721), .Q (n_5605));
  INX1 g41729(.A (n_3439), .Q (n_3438));
  INX1 g41730(.A (n_3437), .Q (instruction[4]));
  NA3I1X2 g41731(.B (n_3422), .C (n_3416), .AN (flush_37507), .Q
       (instruction[0]));
  NA2X4 g41733(.A (n_3429), .B (n_3428), .Q (n_3439));
  AND2X4 g41734(.A (n_3426), .B (n_3420), .Q (n_3437));
  INX1 g41735(.A (instruction[2]), .Q (n_3436));
  INX1 g41737(.A (n_3435), .Q (instruction[18]));
  INX1 g41738(.A (n_3434), .Q (instruction[19]));
  INX1 g41741(.A (instruction[17]), .Q (n_3433));
  BUX4 g41745(.A (n_3431), .Q (\instruction[5]_40139 ));
  INX2 g41746(.A (n_3430), .Q (instruction[3]));
  AO22X1 g41747(.A (n_3287), .B (read_data[11]), .C (n_3285), .D
       (prev_instruction[11]), .Q (\instruction[11]_40800 ));
  AO22X1 g41748(.A (n_3287), .B (read_data[10]), .C (n_3285), .D
       (prev_instruction[10]), .Q (\instruction[10]_39951 ));
  AO22X1 g41749(.A (n_3287), .B (read_data[8]), .C (n_3285), .D
       (prev_instruction[8]), .Q (\instruction[8]_40015 ));
  AO22X1 g41750(.A (n_3287), .B (read_data[9]), .C (n_3285), .D
       (prev_instruction[9]), .Q (\instruction[9]_39983 ));
  AO22X1 g41751(.A (n_3287), .B (read_data[7]), .C (n_3285), .D
       (prev_instruction[7]), .Q (\instruction[7]_39562 ));
  AO22X2 g41754(.A (n_3287), .B (read_data[14]), .C (n_3285), .D
       (prev_instruction[14]), .Q (\instruction[14]_40077 ));
  AO22X1 g41755(.A (n_3394), .B (read_data[2]), .C (n_3393), .D
       (prev_instruction[2]), .Q (instruction[2]));
  AO22X1 g41756(.A (n_3394), .B (read_data[6]), .C (n_3393), .D
       (prev_instruction[6]), .Q (instruction[6]));
  AN22X2 g41757(.A (n_3394), .B (read_data[18]), .C (n_3393), .D
       (prev_instruction[18]), .Q (n_3435));
  AN22X4 g41758(.A (n_3287), .B (read_data[19]), .C (n_3285), .D
       (prev_instruction[19]), .Q (n_3434));
  NA2X4 g41759(.A (n_3421), .B (n_3403), .Q (instruction[17]));
  AO22X2 g41760(.A (n_3287), .B (read_data[5]), .C (n_3285), .D
       (prev_instruction[5]), .Q (n_3431));
  AND2X4 g41761(.A (n_3411), .B (n_3414), .Q (n_3430));
  INX1 g41764(.A (n_3429), .Q (instruction[16]));
  AN21X1 g41767(.A (n_3393), .B (prev_instruction[4]), .C
       (flush_37507), .Q (n_3426));
  NA2I1X4 g41769(.B (n_3402), .AN (n_3397), .Q (instruction[22]));
  AO21X1 g41770(.A (n_3285), .B (prev_instruction[26]), .C (n_3408), .Q
       (instruction[26]));
  AO22X2 g41771(.A (n_3287), .B (read_data[28]), .C (n_3285), .D
       (prev_instruction[28]), .Q (instruction[28]));
  AO22X1 g41772(.A (n_3394), .B (read_data[25]), .C (n_3285), .D
       (prev_instruction[25]), .Q (instruction[25]));
  AO22X2 g41773(.A (n_3394), .B (read_data[29]), .C (n_3285), .D
       (prev_instruction[29]), .Q (instruction[29]));
  AO22X1 g41774(.A (n_3287), .B (read_data[27]), .C (n_3285), .D
       (prev_instruction[27]), .Q (instruction[27]));
  NA2I1X4 g41776(.B (n_3410), .AN (n_3398), .Q (instruction[23]));
  AO22X4 g41777(.A (n_3394), .B (read_data[24]), .C (n_3393), .D
       (prev_instruction[24]), .Q (instruction[24]));
  NO2X4 g41778(.A (n_3400), .B (n_3399), .Q (n_1580));
  NO2X4 g41780(.A (n_3407), .B (n_3406), .Q (n_3429));
  NO2X4 g41781(.A (n_3405), .B (n_3404), .Q (n_3428));
  NA2X1 g41784(.A (n_3393), .B (prev_instruction[0]), .Q (n_3422));
  NA2X1 g41785(.A (n_3393), .B (prev_instruction[17]), .Q (n_3421));
  NA2X1 g41786(.A (n_3394), .B (read_data[4]), .Q (n_3420));
  NA2X1 g41790(.A (n_3394), .B (read_data[0]), .Q (n_3416));
  NA2X1 g41792(.A (n_3394), .B (read_data[3]), .Q (n_3414));
  NA2X1 g41795(.A (n_3393), .B (prev_instruction[3]), .Q (n_3411));
  NA2X2 g41796(.A (n_3392), .B (prev_instruction[23]), .Q (n_3410));
  NO2I1X1 g41797(.B (n_3288), .AN (read_data[13]), .Q (n_3409));
  NO2I1X1 g41798(.B (n_3288), .AN (read_data[26]), .Q (n_3408));
  NO2I1X1 g41799(.B (n_3391), .AN (prev_instruction[16]), .Q (n_3407));
  NO2I1X2 g41800(.B (n_3288), .AN (read_data[16]), .Q (n_3406));
  NO2I1X1 g41801(.B (n_3391), .AN (prev_instruction[15]), .Q (n_3405));
  NO2I1X2 g41802(.B (n_3288), .AN (read_data[15]), .Q (n_3404));
  NA2X1 g41803(.A (n_3394), .B (read_data[17]), .Q (n_3403));
  NA2X2 g41804(.A (n_3392), .B (prev_instruction[22]), .Q (n_3402));
  NO2I1X1 g41806(.B (n_3391), .AN (prev_instruction[21]), .Q (n_3400));
  NO2I1X1 g41807(.B (n_3288), .AN (read_data[21]), .Q (n_3399));
  NO2I1X2 g41808(.B (n_3288), .AN (read_data[23]), .Q (n_3398));
  NO2I1X2 g41809(.B (n_3288), .AN (read_data[22]), .Q (n_3397));
  NO2I1X2 g41810(.B (n_3288), .AN (read_data[20]), .Q (n_3396));
  BUX2 g41817(.A (n_3394), .Q (n_3287));
  NA3I1X4 g41819(.B (n_3389), .C (n_3386), .AN (n_3387), .Q (n_3288));
  AND3X4 g41820(.A (n_3389), .B (n_3388), .C (n_3386), .Q (n_3394));
  BUX4 g41827(.A (n_3393), .Q (n_3285));
  BUX6 g41828(.A (n_3392), .Q (n_3393));
  AND2X4 g41832(.A (n_3390), .B (n_3389), .Q (n_3392));
  NA2X2 g41833(.A (n_3389), .B (n_3390), .Q (n_3391));
  NA2X1 g41834(.A (n_3386), .B (n_3385), .Q (n_6071));
  NA2X4 g41835(.A (n_3386), .B (n_3388), .Q (n_3390));
  INX4 g41836(.A (n_3389), .Q (flush_37507));
  AND3X4 g41837(.A (n_3384), .B (n_3371), .C (current_state[1]), .Q
       (n_3389));
  INX4 g41838(.A (n_3387), .Q (n_3388));
  NA2I1X4 g41839(.B (n_3383), .AN (n_6348), .Q (n_3387));
  NO2X4 g41840(.A (n_3382), .B (halt), .Q (n_3386));
  AND2X1 g41841(.A (n_6348), .B (write_response), .Q
       (store_commit_cycle));
  NA2I1X0 g41842(.B (n_6348), .AN (write_response), .Q (n_3385));
  NO2X2 g41843(.A (current_state[3]), .B (current_state[2]), .Q
       (n_3384));
  NA2X2 g41844(.A (prev_load_request), .B (read_response), .Q (n_3383));
  NO2X2 g41845(.A (n_3363), .B (read_response), .Q (n_3382));
  INX1 g41846(.A (n_5516), .Q (n_3381));
  INX1 g41847(.A (n_5122), .Q (n_3380));
  INX1 g41848(.A (n_5523), .Q (n_3379));
  INX1 g41849(.A (n_4777), .Q (n_3378));
  INX1 g41850(.A (n_5524), .Q (n_3377));
  INX1 g41851(.A (n_5051), .Q (n_3376));
  INX1 g41852(.A (n_5108), .Q (n_3375));
  INX1 g41853(.A (n_4967), .Q (n_3374));
  INX1 g41854(.A (n_4953), .Q (n_3373));
  INX1 g41855(.A (n_4937), .Q (n_3372));
  INX2 g41856(.A (current_state[0]), .Q (n_3371));
  INX1 g41857(.A (n_4963), .Q (n_3370));
  INX1 g41858(.A (n_5515), .Q (n_3369));
  INX1 g41859(.A (n_4882), .Q (n_3368));
  INX1 g41860(.A (n_4776), .Q (n_3367));
  INX1 g41861(.A (n_4646), .Q (n_3366));
  INX1 g41862(.A (n_5115), .Q (n_3365));
  INX1 g41863(.A (n_4962), .Q (n_3364));
  INX1 g41864(.A (n_6347), .Q (n_3363));
  INX1 g41865(.A (n_5457), .Q (n_3362));
  INX1 g41866(.A (n_4938), .Q (n_3361));
  INX1 g41867(.A (n_4881), .Q (n_3360));
  INX1 g41868(.A (n_5512), .Q (n_3359));
  INX1 g41869(.A (n_5397), .Q (n_3358));
  INX1 g41870(.A (n_5116), .Q (n_3357));
  INX1 g41871(.A (n_5396), .Q (n_3356));
  INX1 g41872(.A (n_5456), .Q (n_3355));
  INX1 g41873(.A (n_5050), .Q (n_3354));
  INX1 g41874(.A (n_5513), .Q (n_3353));
  AND2X1 g2(.A (n_3303), .B (n_5150), .Q (n_3283));
  NA2I1X4 g41877(.B (n_3454), .AN (n_3495), .Q (n_3282));
  NA2I1X1 g41878(.B (n_6723), .AN (n_3494), .Q (n_3281));
  NA3I1X1 g41879(.B (n_3436), .C (n_3449), .AN (instruction[6]), .Q
       (n_6598));
  NA2I1X1 g41880(.B (n_3447), .AN (\instruction[5]_40139 ), .Q
       (n_6600));
  AND2X1 g41882(.A (n_176), .B (n_6719), .Q (n_6560));
  INX1 g41884(.A (n_3298), .Q (n_3297));
  INX1 g41886(.A (n_3301), .Q (n_3300));
  INX1 g41892(.A (n_3305), .Q (n_3304));
  AND2X1 g41894(.A (n_3973), .B (n_3989), .Q (n_3325));
  AND2X1 g41898(.A (n_3978), .B (n_3763), .Q (n_3329));
  AND2X1 g41900(.A (n_3981), .B (n_3997), .Q (n_3326));
  AND2X1 g41910(.A (n_3942), .B (n_3943), .Q (n_3323));
  AND2X1 g41912(.A (n_3975), .B (n_3991), .Q (n_3324));
  AND2X1 g41914(.A (n_3976), .B (n_3992), .Q (n_3328));
  AND2X1 g41916(.A (n_3938), .B (n_3939), .Q (n_3322));
  AO221X1 g41918(.A (n_5266), .B (n_3520), .C (n_3518), .D (n_5272), .E
       (n_3703), .Q (n_3315));
  AND6X1 g41920(.A (n_4352), .B (n_4268), .C (n_4140), .D (n_4149), .E
       (n_4150), .F (n_4141), .Q (n_3352));
  AND2X1 g41922(.A (n_3816), .B (n_3817), .Q (n_3316));
  AND2X1 g41924(.A (n_3810), .B (n_3811), .Q (n_3311));
  AND2X1 g41930(.A (n_3915), .B (n_3955), .Q (n_3321));
  AND2X1 g41932(.A (n_3913), .B (n_3953), .Q (n_3317));
  AND2X1 g41936(.A (n_3908), .B (n_3948), .Q (n_3318));
  AND2X1 g41938(.A (n_3820), .B (n_3828), .Q (n_3310));
  AND2X1 g41940(.A (n_3819), .B (n_3827), .Q (n_3309));
  AND6X1 g41942(.A (n_6644), .B (n_4267), .C (n_4138), .D (n_4145), .E
       (n_4137), .F (n_4146), .Q (n_3351));
  AND6X1 g41944(.A (n_4314), .B (n_4315), .C (n_4037), .D (n_4039), .E
       (n_4049), .F (n_4051), .Q (n_3337));
  AND6X1 g41946(.A (n_4329), .B (n_4328), .C (n_4115), .D (n_4084), .E
       (n_4086), .F (n_4085), .Q (n_3347));
  AND6X1 g41948(.A (n_4355), .B (n_4356), .C (n_4184), .D (n_4189), .E
       (n_4190), .F (n_4191), .Q (n_3339));
  AND6X1 g41950(.A (n_4064), .B (n_4284), .C (n_4009), .D (n_4242), .E
       (n_3905), .F (n_3945), .Q (n_3331));
  AND6X1 g41952(.A (n_3324), .B (n_3328), .C (n_3977), .D (n_3974), .E
       (n_3990), .F (n_3993), .Q (n_3333));
  AND6X1 g41954(.A (n_6646), .B (n_4265), .C (n_4108), .D (n_4107), .E
       (n_4078), .F (n_4079), .Q (n_3342));
  AND2X2 g41956(.A (n_3499), .B (n_3484), .Q (n_3303));
  AND6X1 g41958(.A (n_6650), .B (n_4165), .C (n_4258), .D (n_4118), .E
       (n_4117), .F (n_4119), .Q (n_3346));
  AND6X1 g41960(.A (n_4280), .B (n_4275), .C (n_4194), .D (n_4195), .E
       (n_3980), .F (n_4188), .Q (n_3336));
  AND6X1 g41962(.A (n_4283), .B (n_3323), .C (n_4063), .D (n_4008), .E
       (n_4006), .F (n_4007), .Q (n_3332));
  AND6X1 g41964(.A (n_6647), .B (n_4161), .C (n_6660), .D (n_4160), .E
       (n_4109), .F (n_4080), .Q (n_3343));
  AND6X1 g41966(.A (n_6645), .B (n_4266), .C (n_4111), .D (n_4082), .E
       (n_4083), .F (n_4112), .Q (n_3344));
  AND6X1 g41968(.A (n_4358), .B (n_4338), .C (n_4176), .D (n_4175), .E
       (n_4147), .F (n_4148), .Q (n_3349));
  AND6X1 g41970(.A (n_6656), .B (n_6778), .C (n_3982), .D (n_3998), .E
       (n_3983), .F (n_3999), .Q (n_3335));
  AND6X1 g41972(.A (n_6776), .B (n_4331), .C (n_4172), .D (n_4171), .E
       (n_4142), .F (n_4151), .Q (n_3350));
  AND6X1 g41974(.A (n_6777), .B (n_4179), .C (n_4153), .D (n_4152), .E
       (n_4154), .F (n_4264), .Q (n_3348));
  AND6X1 g41976(.A (n_4344), .B (n_4168), .C (n_4317), .D (n_4124), .E
       (n_4055), .F (n_4056), .Q (n_3340));
  AND6X1 g41978(.A (n_6649), .B (n_4259), .C (n_4048), .D (n_4046), .E
       (n_4058), .F (n_4060), .Q (n_3338));
  AND6X1 g41980(.A (n_6654), .B (n_4130), .C (n_4092), .D (n_4090), .E
       (n_4091), .F (n_4250), .Q (n_3341));
  AND6X1 g41982(.A (n_6643), .B (n_4156), .C (n_6659), .D (n_4155), .E
       (n_4105), .F (n_4076), .Q (n_3345));
  AND6X1 g41984(.A (n_6652), .B (n_6697), .C (n_3984), .D (n_4000), .E
       (n_3985), .F (n_4001), .Q (n_3334));
  INX2 g41986(.A (n_3428), .Q (instruction[15]));
  AND2X1 g41988(.A (n_5605), .B (\instruction[14]_40077 ), .Q (n_6457));
  INX2 g41990(.A (n_3489), .Q (n_3293));
  INX2 g41992(.A (n_3488), .Q (n_3292));
  INX1 g41995(.A (n_3296), .Q (n_3294));
  DFRQX1 \csr_mepc_reg[0] (.C (rc_gclk_205556), .D (n_3233), .Q
       (n_3260));
  DFRQX1 \csr_mepc_reg[1] (.C (rc_gclk_205556), .D (n_3234), .Q
       (n_3261));
  DFRQX1 csr_mip_meip_reg(.C (clock), .D (n_1781), .Q (n_3262));
  DFRQX1 \csr_mip_mfip_reg[0] (.C (clock), .D (n_1791), .Q (n_3265));
  DFRQX1 \csr_mip_mfip_reg[10] (.C (clock), .D (n_1795), .Q (n_3275));
  DFRQX1 \csr_mip_mfip_reg[11] (.C (clock), .D (n_1792), .Q (n_3276));
  DFRQX1 \csr_mip_mfip_reg[12] (.C (clock), .D (n_1783), .Q (n_3277));
  DFRQX1 \csr_mip_mfip_reg[13] (.C (clock), .D (n_1788), .Q (n_3278));
  DFRQX1 \csr_mip_mfip_reg[14] (.C (clock), .D (n_1789), .Q (n_3279));
  DFRQX1 \csr_mip_mfip_reg[15] (.C (clock), .D (n_1787), .Q (n_3280));
  DFRQX1 \csr_mip_mfip_reg[1] (.C (clock), .D (n_1780), .Q (n_3266));
  DFRQX1 \csr_mip_mfip_reg[2] (.C (clock), .D (n_1793), .Q (n_3267));
  DFRQX1 \csr_mip_mfip_reg[3] (.C (clock), .D (n_1779), .Q (n_3268));
  DFRQX1 \csr_mip_mfip_reg[4] (.C (clock), .D (n_1786), .Q (n_3269));
  DFRQX1 \csr_mip_mfip_reg[5] (.C (clock), .D (n_1778), .Q (n_3270));
  DFRQX1 \csr_mip_mfip_reg[6] (.C (clock), .D (n_1784), .Q (n_3271));
  DFRQX1 \csr_mip_mfip_reg[7] (.C (clock), .D (n_1785), .Q (n_3272));
  DFRQX1 \csr_mip_mfip_reg[8] (.C (clock), .D (n_1794), .Q (n_3273));
  DFRQX1 \csr_mip_mfip_reg[9] (.C (clock), .D (n_1777), .Q (n_3274));
  DFRQX1 csr_mip_msip_reg(.C (clock), .D (n_1790), .Q (n_3264));
  DFRQX1 csr_mip_mtip_reg(.C (clock), .D (n_1782), .Q (n_3263));
  DFRQX1 \csr_utime_reg[0] (.C (clock), .D (real_time_clock[0]), .Q
       (csr_utime[0]));
  DFRQX1 \csr_utime_reg[10] (.C (clock), .D (real_time_clock[10]), .Q
       (csr_utime[10]));
  DFRQX1 \csr_utime_reg[11] (.C (clock), .D (real_time_clock[11]), .Q
       (csr_utime[11]));
  DFRQX1 \csr_utime_reg[12] (.C (clock), .D (real_time_clock[12]), .Q
       (csr_utime[12]));
  DFRQX1 \csr_utime_reg[13] (.C (clock), .D (real_time_clock[13]), .Q
       (csr_utime[13]));
  DFRQX1 \csr_utime_reg[14] (.C (clock), .D (real_time_clock[14]), .Q
       (csr_utime[14]));
  DFRQX1 \csr_utime_reg[15] (.C (clock), .D (real_time_clock[15]), .Q
       (csr_utime[15]));
  DFRQX1 \csr_utime_reg[16] (.C (clock), .D (real_time_clock[16]), .Q
       (csr_utime[16]));
  DFRQX1 \csr_utime_reg[17] (.C (clock), .D (real_time_clock[17]), .Q
       (csr_utime[17]));
  DFRQX1 \csr_utime_reg[18] (.C (clock), .D (real_time_clock[18]), .Q
       (csr_utime[18]));
  DFRQX1 \csr_utime_reg[19] (.C (clock), .D (real_time_clock[19]), .Q
       (csr_utime[19]));
  DFRQX1 \csr_utime_reg[1] (.C (clock), .D (real_time_clock[1]), .Q
       (csr_utime[1]));
  DFRQX1 \csr_utime_reg[20] (.C (clock), .D (real_time_clock[20]), .Q
       (csr_utime[20]));
  DFRQX1 \csr_utime_reg[21] (.C (clock), .D (real_time_clock[21]), .Q
       (csr_utime[21]));
  DFRQX1 \csr_utime_reg[22] (.C (clock), .D (real_time_clock[22]), .Q
       (csr_utime[22]));
  DFRQX1 \csr_utime_reg[23] (.C (clock), .D (real_time_clock[23]), .Q
       (csr_utime[23]));
  DFRQX1 \csr_utime_reg[24] (.C (clock), .D (real_time_clock[24]), .Q
       (csr_utime[24]));
  DFRQX1 \csr_utime_reg[25] (.C (clock), .D (real_time_clock[25]), .Q
       (csr_utime[25]));
  DFRQX1 \csr_utime_reg[26] (.C (clock), .D (real_time_clock[26]), .Q
       (csr_utime[26]));
  DFRQX1 \csr_utime_reg[27] (.C (clock), .D (real_time_clock[27]), .Q
       (csr_utime[27]));
  DFRQX1 \csr_utime_reg[28] (.C (clock), .D (real_time_clock[28]), .Q
       (csr_utime[28]));
  DFRQX1 \csr_utime_reg[29] (.C (clock), .D (real_time_clock[29]), .Q
       (csr_utime[29]));
  DFRQX1 \csr_utime_reg[2] (.C (clock), .D (real_time_clock[2]), .Q
       (csr_utime[2]));
  DFRQX1 \csr_utime_reg[30] (.C (clock), .D (real_time_clock[30]), .Q
       (csr_utime[30]));
  DFRQX1 \csr_utime_reg[31] (.C (clock), .D (real_time_clock[31]), .Q
       (csr_utime[31]));
  DFRQX1 \csr_utime_reg[32] (.C (clock), .D (real_time_clock[32]), .Q
       (csr_utime[32]));
  DFRQX1 \csr_utime_reg[33] (.C (clock), .D (real_time_clock[33]), .Q
       (csr_utime[33]));
  DFRQX1 \csr_utime_reg[34] (.C (clock), .D (real_time_clock[34]), .Q
       (csr_utime[34]));
  DFRQX1 \csr_utime_reg[35] (.C (clock), .D (real_time_clock[35]), .Q
       (csr_utime[35]));
  DFRQX1 \csr_utime_reg[36] (.C (clock), .D (real_time_clock[36]), .Q
       (csr_utime[36]));
  DFRQX1 \csr_utime_reg[37] (.C (clock), .D (real_time_clock[37]), .Q
       (csr_utime[37]));
  DFRQX1 \csr_utime_reg[38] (.C (clock), .D (real_time_clock[38]), .Q
       (csr_utime[38]));
  DFRQX1 \csr_utime_reg[39] (.C (clock), .D (real_time_clock[39]), .Q
       (csr_utime[39]));
  DFRQX1 \csr_utime_reg[3] (.C (clock), .D (real_time_clock[3]), .Q
       (csr_utime[3]));
  DFRQX1 \csr_utime_reg[40] (.C (clock), .D (real_time_clock[40]), .Q
       (csr_utime[40]));
  DFRQX1 \csr_utime_reg[41] (.C (clock), .D (real_time_clock[41]), .Q
       (csr_utime[41]));
  DFRQX1 \csr_utime_reg[42] (.C (clock), .D (real_time_clock[42]), .Q
       (csr_utime[42]));
  DFRQX1 \csr_utime_reg[43] (.C (clock), .D (real_time_clock[43]), .Q
       (csr_utime[43]));
  DFRQX1 \csr_utime_reg[44] (.C (clock), .D (real_time_clock[44]), .Q
       (csr_utime[44]));
  DFRQX1 \csr_utime_reg[45] (.C (clock), .D (real_time_clock[45]), .Q
       (csr_utime[45]));
  DFRQX1 \csr_utime_reg[46] (.C (clock), .D (real_time_clock[46]), .Q
       (csr_utime[46]));
  DFRQX1 \csr_utime_reg[47] (.C (clock), .D (real_time_clock[47]), .Q
       (csr_utime[47]));
  DFRQX1 \csr_utime_reg[48] (.C (clock), .D (real_time_clock[48]), .Q
       (csr_utime[48]));
  DFRQX1 \csr_utime_reg[49] (.C (clock), .D (real_time_clock[49]), .Q
       (csr_utime[49]));
  DFRQX1 \csr_utime_reg[4] (.C (clock), .D (real_time_clock[4]), .Q
       (csr_utime[4]));
  DFRQX1 \csr_utime_reg[50] (.C (clock), .D (real_time_clock[50]), .Q
       (csr_utime[50]));
  DFRQX1 \csr_utime_reg[51] (.C (clock), .D (real_time_clock[51]), .Q
       (csr_utime[51]));
  DFRQX1 \csr_utime_reg[52] (.C (clock), .D (real_time_clock[52]), .Q
       (csr_utime[52]));
  DFRQX1 \csr_utime_reg[53] (.C (clock), .D (real_time_clock[53]), .Q
       (csr_utime[53]));
  DFRQX1 \csr_utime_reg[54] (.C (clock), .D (real_time_clock[54]), .Q
       (csr_utime[54]));
  DFRQX1 \csr_utime_reg[55] (.C (clock), .D (real_time_clock[55]), .Q
       (csr_utime[55]));
  DFRQX1 \csr_utime_reg[56] (.C (clock), .D (real_time_clock[56]), .Q
       (csr_utime[56]));
  DFRQX1 \csr_utime_reg[57] (.C (clock), .D (real_time_clock[57]), .Q
       (csr_utime[57]));
  DFRQX1 \csr_utime_reg[58] (.C (clock), .D (real_time_clock[58]), .Q
       (csr_utime[58]));
  DFRQX1 \csr_utime_reg[59] (.C (clock), .D (real_time_clock[59]), .Q
       (csr_utime[59]));
  DFRQX1 \csr_utime_reg[5] (.C (clock), .D (real_time_clock[5]), .Q
       (csr_utime[5]));
  DFRQX1 \csr_utime_reg[60] (.C (clock), .D (real_time_clock[60]), .Q
       (csr_utime[60]));
  DFRQX1 \csr_utime_reg[61] (.C (clock), .D (real_time_clock[61]), .Q
       (csr_utime[61]));
  DFRQX1 \csr_utime_reg[62] (.C (clock), .D (real_time_clock[62]), .Q
       (csr_utime[62]));
  DFRQX1 \csr_utime_reg[63] (.C (clock), .D (real_time_clock[63]), .Q
       (csr_utime[63]));
  DFRQX1 \csr_utime_reg[6] (.C (clock), .D (real_time_clock[6]), .Q
       (csr_utime[6]));
  DFRQX1 \csr_utime_reg[7] (.C (clock), .D (real_time_clock[7]), .Q
       (csr_utime[7]));
  DFRQX1 \csr_utime_reg[8] (.C (clock), .D (real_time_clock[8]), .Q
       (csr_utime[8]));
  DFRQX1 \csr_utime_reg[9] (.C (clock), .D (real_time_clock[9]), .Q
       (csr_utime[9]));
  DFRQX1 reset_reg_reg(.C (clock), .D (reset), .Q (reset_reg));
  AO211X1 g61576(.A (n_3256), .B (n_6238), .C (n_6506), .D (n_3257), .Q
       (n_5627));
  NA2X4 g61577(.A (n_3258), .B (n_1809), .Q (n_4534));
  AO22X2 g61579(.A (instruction_address[0]), .B (n_1663), .C (n_1585),
       .D (prev_rw_address[0]), .Q (rw_address[0]));
  AO22X2 g61580(.A (n_1663), .B (instruction_address[1]), .C (n_1585),
       .D (prev_rw_address[1]), .Q (rw_address[1]));
  NA2X2 g61582(.A (n_1902), .B (csr_data_out[0]), .Q (n_3258));
  OR5X1 g61583(.A (n_6508), .B (n_6507), .C (n_6515), .D (n_6517), .E
       (n_6520), .Q (n_3257));
  NA6I3X1 g61584(.D (n_1577), .E (n_3239), .F (n_3237), .AN (n_3252),
       .BN (n_3244), .CN (n_1572), .Q (n_3256));
  NA3X1 g61585(.A (n_2140), .B (n_3253), .C (n_2024), .Q
       (csr_data_out[0]));
  NA3X1 g61586(.A (n_3255), .B (n_2124), .C (n_2122), .Q
       (csr_data_out[1]));
  NO3X1 g61587(.A (n_3254), .B (n_1982), .C (n_1922), .Q (n_6503));
  NO2X1 g61588(.A (n_3254), .B (n_1930), .Q (n_6505));
  NO2X1 g61589(.A (n_3254), .B (n_1921), .Q (n_6506));
  NO2X1 g61590(.A (n_3254), .B (n_1926), .Q (n_6504));
  AN221X1 g61591(.A (csr_minstret[1]), .B (n_6625), .C
       (csr_mcycle[33]), .D (n_1937), .E (n_3251), .Q (n_3255));
  AO22X1 g61592(.A (n_6529), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[1]), .Q (instruction_address[1]));
  AO22X1 g61593(.A (n_6528), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[0]), .Q (instruction_address[0]));
  NO3X1 g61594(.A (n_3250), .B (n_1664), .C (n_1920), .Q (n_6508));
  NO2X1 g61595(.A (n_3250), .B (n_1984), .Q (n_6507));
  NA3X1 g61596(.A (n_3249), .B (n_1984), .C (n_5542), .Q (n_3254));
  AN221X1 g61597(.A (csr_mcause[0]), .B (n_2012), .C (csr_mtval[0]), .D
       (n_2016), .E (n_3248), .Q (n_3253));
  NO2X1 g61598(.A (n_1577), .B (n_1723), .Q (n_6509));
  NA3X1 g61599(.A (n_3247), .B (n_3245), .C (n_3246), .Q (n_3252));
  AO222X1 g61600(.A (n_3261), .B (n_2014), .C (csr_minstret[33]), .D
       (n_1938), .E (csr_mscratch[1]), .F (n_1970), .Q (n_3251));
  NO2X1 g61601(.A (n_3247), .B (n_1723), .Q (n_6512));
  AO22X2 g61602(.A (write_request), .B (n_2792), .C (n_1585), .D
       (prev_write_strobe[3]), .Q (write_strobe[3]));
  AO22X2 g61603(.A (write_request), .B (n_2959), .C (n_1585), .D
       (prev_write_strobe[2]), .Q (write_strobe[2]));
  AO22X2 g61604(.A (write_request), .B (n_2691), .C (n_1585), .D
       (prev_write_strobe[1]), .Q (write_strobe[1]));
  AND2X1 g61605(.A (n_1572), .B (n_6238), .Q (n_6514));
  AND2X1 g61606(.A (n_3244), .B (n_6238), .Q (n_6513));
  AO22X2 g61607(.A (write_request), .B (n_2795), .C (n_1585), .D
       (prev_write_strobe[0]), .Q (write_strobe[0]));
  INX1 g61608(.A (n_3249), .Q (n_3250));
  AO22X1 g61609(.A (n_2014), .B (n_3260), .C (n_1970), .D
       (csr_mscratch[0]), .Q (n_3248));
  NO2X1 g61610(.A (n_3246), .B (n_1723), .Q (n_6511));
  NO2X1 g61611(.A (n_3245), .B (n_1723), .Q (n_6510));
  ON21X1 g61612(.A (n_3225), .B (n_1848), .C (n_3243), .Q (n_6529));
  AO22X1 g61613(.A (n_211), .B (n_3260), .C (n_3223), .D
       (program_counter[0]), .Q (n_6528));
  NO3X1 g61615(.A (n_1574), .B (n_1723), .C (n_1985), .Q (n_3249));
  AO222X2 g61616(.A (instruction_address[30]), .B (n_1663), .C
       (n_5704), .D (n_3230), .E (prev_rw_address[30]), .F (n_1585), .Q
       (rw_address[30]));
  AO222X2 g61617(.A (instruction_address[8]), .B (n_1663), .C (n_5709),
       .D (n_3230), .E (prev_rw_address[8]), .F (n_1585), .Q
       (rw_address[8]));
  AO222X2 g61618(.A (instruction_address[4]), .B (n_1663), .C (n_5713),
       .D (n_3230), .E (prev_rw_address[4]), .F (n_1585), .Q
       (rw_address[4]));
  AO222X2 g61619(.A (instruction_address[7]), .B (n_1663), .C (n_5710),
       .D (n_3230), .E (prev_rw_address[7]), .F (n_1585), .Q
       (rw_address[7]));
  AO222X2 g61620(.A (instruction_address[2]), .B (n_1663), .C (n_5716),
       .D (n_3230), .E (prev_rw_address[2]), .F (n_1585), .Q
       (rw_address[2]));
  AO222X2 g61621(.A (instruction_address[6]), .B (n_1663), .C (n_5711),
       .D (n_3230), .E (prev_rw_address[6]), .F (n_1585), .Q
       (rw_address[6]));
  AO222X2 g61622(.A (instruction_address[5]), .B (n_1663), .C (n_5712),
       .D (n_3230), .E (prev_rw_address[5]), .F (n_1585), .Q
       (rw_address[5]));
  AO222X2 g61623(.A (instruction_address[3]), .B (n_1663), .C (n_5714),
       .D (n_3230), .E (prev_rw_address[3]), .F (n_1585), .Q
       (rw_address[3]));
  AO222X2 g61624(.A (instruction_address[31]), .B (n_1663), .C
       (n_5682), .D (n_3230), .E (prev_rw_address[31]), .F (n_1585), .Q
       (rw_address[31]));
  AO222X2 g61625(.A (instruction_address[9]), .B (n_1663), .C (n_5708),
       .D (n_3230), .E (prev_rw_address[9]), .F (n_1585), .Q
       (rw_address[9]));
  AO222X2 g61626(.A (instruction_address[29]), .B (n_1663), .C
       (n_5715), .D (n_3230), .E (prev_rw_address[29]), .F (n_1585), .Q
       (rw_address[29]));
  AO222X2 g61627(.A (instruction_address[28]), .B (n_1663), .C
       (n_5717), .D (n_3230), .E (prev_rw_address[28]), .F (n_1585), .Q
       (rw_address[28]));
  AO222X2 g61628(.A (instruction_address[27]), .B (n_1663), .C
       (n_5718), .D (n_3230), .E (prev_rw_address[27]), .F (n_1585), .Q
       (rw_address[27]));
  AO222X2 g61629(.A (instruction_address[26]), .B (n_1663), .C
       (n_5719), .D (n_3230), .E (prev_rw_address[26]), .F (n_1585), .Q
       (rw_address[26]));
  AO222X2 g61630(.A (instruction_address[25]), .B (n_1663), .C
       (n_5720), .D (n_3230), .E (prev_rw_address[25]), .F (n_1585), .Q
       (rw_address[25]));
  AO222X2 g61631(.A (instruction_address[24]), .B (n_1663), .C
       (n_5721), .D (n_3230), .E (prev_rw_address[24]), .F (n_1585), .Q
       (rw_address[24]));
  AO222X2 g61632(.A (instruction_address[23]), .B (n_1663), .C
       (n_5722), .D (n_3230), .E (prev_rw_address[23]), .F (n_1585), .Q
       (rw_address[23]));
  AO222X2 g61633(.A (instruction_address[22]), .B (n_1663), .C
       (n_5684), .D (n_3230), .E (prev_rw_address[22]), .F (n_1585), .Q
       (rw_address[22]));
  AO222X2 g61634(.A (instruction_address[21]), .B (n_1663), .C
       (n_5686), .D (n_3230), .E (prev_rw_address[21]), .F (n_1585), .Q
       (rw_address[21]));
  AO222X2 g61636(.A (instruction_address[11]), .B (n_1663), .C
       (n_5706), .D (n_3230), .E (prev_rw_address[11]), .F (n_1585), .Q
       (rw_address[11]));
  AO222X2 g61637(.A (instruction_address[19]), .B (n_1663), .C
       (n_5690), .D (n_3230), .E (prev_rw_address[19]), .F (n_1585), .Q
       (rw_address[19]));
  AO222X2 g61638(.A (instruction_address[18]), .B (n_1663), .C
       (n_5692), .D (n_3230), .E (prev_rw_address[18]), .F (n_1585), .Q
       (rw_address[18]));
  AO222X2 g61639(.A (instruction_address[17]), .B (n_1663), .C
       (n_5694), .D (n_3230), .E (prev_rw_address[17]), .F (n_1585), .Q
       (rw_address[17]));
  AO222X2 g61640(.A (instruction_address[16]), .B (n_1663), .C
       (n_5696), .D (n_3230), .E (prev_rw_address[16]), .F (n_1585), .Q
       (rw_address[16]));
  AO222X2 g61641(.A (instruction_address[15]), .B (n_1663), .C
       (n_5698), .D (n_3230), .E (prev_rw_address[15]), .F (n_1585), .Q
       (rw_address[15]));
  AO222X2 g61642(.A (instruction_address[14]), .B (n_1663), .C
       (n_5700), .D (n_3230), .E (prev_rw_address[14]), .F (n_1585), .Q
       (rw_address[14]));
  AO222X2 g61643(.A (instruction_address[13]), .B (n_1663), .C
       (n_5702), .D (n_3230), .E (prev_rw_address[13]), .F (n_1585), .Q
       (rw_address[13]));
  AO222X2 g61644(.A (instruction_address[12]), .B (n_1663), .C
       (n_5705), .D (n_3230), .E (prev_rw_address[12]), .F (n_1585), .Q
       (rw_address[12]));
  AO222X2 g61645(.A (instruction_address[20]), .B (n_1663), .C
       (n_5688), .D (n_3230), .E (prev_rw_address[20]), .F (n_1585), .Q
       (rw_address[20]));
  AO222X2 g61646(.A (instruction_address[10]), .B (n_1663), .C
       (n_5707), .D (n_3230), .E (prev_rw_address[10]), .F (n_1585), .Q
       (rw_address[10]));
  NA2X1 g61647(.A (n_211), .B (n_3261), .Q (n_3243));
  NO3X1 g61648(.A (n_3240), .B (n_1723), .C (n_1912), .Q (n_6515));
  OR4X1 g61649(.A (n_3240), .B (n_1980), .C (n_1911), .D (n_1924), .Q
       (n_3247));
  NA2X1 g61651(.A (n_3242), .B (n_1975), .Q (n_3246));
  OR4X1 g61652(.A (n_3241), .B (n_1975), .C (n_1664), .D (n_1917), .Q
       (n_3245));
  NO3X1 g61654(.A (n_3240), .B (n_1980), .C (n_1910), .Q (n_3244));
  INX1 g61655(.A (n_3241), .Q (n_3242));
  AO22X1 g61656(.A (n_3232), .B (n_1799), .C (n_1585), .D (n_6347), .Q
       (read_request));
  AN211X1 g61657(.A (n_3228), .B (n_1983), .C (n_3226), .D (n_3236), .Q
       (n_3239));
  NA2X1 g61659(.A (n_3238), .B (n_2086), .Q (n_3241));
  NA2X1 g61660(.A (n_3238), .B (n_5542), .Q (n_3240));
  AND2X1 g61661(.A (n_3236), .B (n_6238), .Q (n_6516));
  ON21X1 g61662(.A (n_2015), .B (n_1565), .C (n_3235), .Q (n_6499));
  ON21X1 g61663(.A (n_2013), .B (n_1565), .C (n_3235), .Q (n_6479));
  AO22X2 g61666(.A (n_3231), .B (n_1799), .C (n_1585), .D (n_6348), .Q
       (write_request));
  AO22X1 g61667(.A (n_6537), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[8]), .Q (instruction_address[8]));
  AO22X1 g61668(.A (n_6536), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[7]), .Q (instruction_address[7]));
  AO22X1 g61669(.A (n_6534), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[5]), .Q (instruction_address[5]));
  AO22X1 g61670(.A (n_6527), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[28]), .Q (instruction_address[28]));
  AO22X1 g61671(.A (n_6546), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[16]), .Q (instruction_address[16]));
  AO22X1 g61672(.A (n_6544), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[14]), .Q (instruction_address[14]));
  AO22X1 g61673(.A (n_6541), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[12]), .Q (instruction_address[12]));
  AO22X1 g61674(.A (n_6540), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[11]), .Q (instruction_address[11]));
  AO22X1 g61675(.A (n_6539), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[10]), .Q (instruction_address[10]));
  AO22X1 g61676(.A (n_6538), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[9]), .Q (instruction_address[9]));
  AO22X1 g61677(.A (n_6535), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[6]), .Q (instruction_address[6]));
  AO22X1 g61678(.A (n_6533), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[4]), .Q (instruction_address[4]));
  AO22X1 g61679(.A (n_6532), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[3]), .Q (instruction_address[3]));
  AO22X1 g61680(.A (n_6553), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[31]), .Q (instruction_address[31]));
  AO22X1 g61681(.A (n_6542), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[30]), .Q (instruction_address[30]));
  AO22X1 g61682(.A (n_6531), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[29]), .Q (instruction_address[29]));
  AO22X1 g61683(.A (n_6526), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[27]), .Q (instruction_address[27]));
  AO22X1 g61684(.A (n_6525), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[26]), .Q (instruction_address[26]));
  AO22X1 g61685(.A (n_6524), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[25]), .Q (instruction_address[25]));
  ON21X1 g61686(.A (n_1661), .B (n_1723), .C (n_121), .Q (n_5628));
  AND3X1 g61687(.A (take_trap_39145), .B (program_counter[1]), .C
       (n_121), .Q (n_3234));
  AND3X1 g61688(.A (take_trap_39145), .B (program_counter[0]), .C
       (n_121), .Q (n_3233));
  AO22X1 g61689(.A (n_6551), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[21]), .Q (instruction_address[21]));
  AO22X1 g61690(.A (n_6550), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[20]), .Q (instruction_address[20]));
  AO22X1 g61691(.A (n_6549), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[19]), .Q (instruction_address[19]));
  AO22X1 g61692(.A (n_6548), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[18]), .Q (instruction_address[18]));
  AO22X1 g61693(.A (n_6547), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[17]), .Q (instruction_address[17]));
  AO22X1 g61694(.A (n_6545), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[15]), .Q (instruction_address[15]));
  AO22X1 g61695(.A (n_6543), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[13]), .Q (instruction_address[13]));
  AO22X1 g61696(.A (n_6530), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[2]), .Q (instruction_address[2]));
  AND4X1 g61697(.A (n_3229), .B (n_1979), .C (n_1973), .D (n_1913), .Q
       (n_3238));
  AND4X1 g61698(.A (n_3229), .B (n_6238), .C (n_1979), .D (n_1972), .Q
       (n_6517));
  NA2X1 g61699(.A (n_3229), .B (n_1978), .Q (n_3237));
  AND5X1 g61700(.A (n_3229), .B (n_1973), .C (n_1914), .D (n_5542), .E
       (n_1909), .Q (n_3236));
  AN21X1 g61701(.A (n_1662), .B (n_1688), .C (n_1748), .Q (n_3235));
  AO22X1 g61702(.A (n_6523), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[24]), .Q (instruction_address[24]));
  AO22X1 g61703(.A (n_6522), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[23]), .Q (instruction_address[23]));
  AO22X1 g61704(.A (n_6552), .B (n_1722), .C (n_1721), .D
       (prev_instruction_address[22]), .Q (instruction_address[22]));
  INX1 g61706(.A (n_3231), .Q (n_3232));
  NO2X1 g61707(.A (n_1662), .B (n_1823), .Q (n_3231));
  AND3X1 g61708(.A (n_1661), .B (n_2085), .C (n_1799), .Q (n_3230));
  NA2X1 g61709(.A (n_1661), .B (n_1974), .Q (load_request_BAR));
  AND2X1 g61710(.A (n_3226), .B (n_6238), .Q (n_6519));
  NO2X1 g61711(.A (n_3227), .B (n_1983), .Q (n_3229));
  AO221X1 g61712(.A (n_5579), .B (n_3223), .C (n_5710), .D (n_3220), .E
       (n_1959), .Q (n_6536));
  AO221X1 g61713(.A (n_5578), .B (n_3223), .C (n_5711), .D (n_3220), .E
       (n_1958), .Q (n_6535));
  AO221X1 g61714(.A (n_5603), .B (n_3223), .C (n_5682), .D (n_3220), .E
       (n_2000), .Q (n_6553));
  AO221X1 g61715(.A (n_5602), .B (n_3223), .C (n_5704), .D (n_3220), .E
       (n_1999), .Q (n_6542));
  AO221X1 g61716(.A (n_5599), .B (n_3223), .C (n_5718), .D (n_3220), .E
       (n_2005), .Q (n_6526));
  AO221X1 g61717(.A (n_5596), .B (n_3223), .C (n_5721), .D (n_3220), .E
       (n_1989), .Q (n_6523));
  AO221X1 g61718(.A (n_5595), .B (n_3223), .C (n_5722), .D (n_3220), .E
       (n_2004), .Q (n_6522));
  AO221X1 g61719(.A (n_5592), .B (n_3223), .C (n_5688), .D (n_3220), .E
       (n_1988), .Q (n_6550));
  AO221X1 g61720(.A (n_5591), .B (n_3223), .C (n_5690), .D (n_3220), .E
       (n_2003), .Q (n_6549));
  AO221X1 g61721(.A (n_5589), .B (n_3223), .C (n_5694), .D (n_3220), .E
       (n_1987), .Q (n_6547));
  AO221X1 g61722(.A (n_5582), .B (n_3223), .C (n_5707), .D (n_3220), .E
       (n_1965), .Q (n_6539));
  AO221X1 g61723(.A (n_5581), .B (n_3223), .C (n_5708), .D (n_3220), .E
       (n_1962), .Q (n_6538));
  AO221X1 g61724(.A (n_5580), .B (n_3223), .C (n_5709), .D (n_3220), .E
       (n_1960), .Q (n_6537));
  AO221X1 g61725(.A (n_5577), .B (n_3223), .C (n_5712), .D (n_3220), .E
       (n_1957), .Q (n_6534));
  AO221X1 g61726(.A (n_5576), .B (n_3223), .C (n_5713), .D (n_3220), .E
       (n_1956), .Q (n_6533));
  AO221X1 g61727(.A (n_5575), .B (n_3223), .C (n_5714), .D (n_3220), .E
       (n_1955), .Q (n_6532));
  ON221X1 g61728(.A (program_counter[2]), .B (n_3222), .C (n_2118), .D
       (n_3221), .E (n_1963), .Q (n_6530));
  INX1 g61729(.A (n_3227), .Q (n_3228));
  INX1 g61738(.A (n_1662), .Q (n_1661));
  AO221X1 g61739(.A (n_5601), .B (n_3223), .C (n_5715), .D (n_3220), .E
       (n_1998), .Q (n_6531));
  AO221X1 g61740(.A (n_5600), .B (n_3223), .C (n_5717), .D (n_3220), .E
       (n_1991), .Q (n_6527));
  AO221X1 g61741(.A (n_5598), .B (n_3223), .C (n_5719), .D (n_3220), .E
       (n_2009), .Q (n_6525));
  AO221X1 g61742(.A (n_5597), .B (n_3223), .C (n_5720), .D (n_3220), .E
       (n_1996), .Q (n_6524));
  AO221X1 g61743(.A (n_5594), .B (n_3223), .C (n_5684), .D (n_3220), .E
       (n_1995), .Q (n_6552));
  AO221X1 g61744(.A (n_5593), .B (n_3223), .C (n_5686), .D (n_3220), .E
       (n_1994), .Q (n_6551));
  AO221X1 g61745(.A (n_5590), .B (n_3223), .C (n_5692), .D (n_3220), .E
       (n_1993), .Q (n_6548));
  AO221X1 g61746(.A (n_5588), .B (n_3223), .C (n_5696), .D (n_3220), .E
       (n_1966), .Q (n_6546));
  AO221X1 g61747(.A (n_5587), .B (n_3223), .C (n_5698), .D (n_3220), .E
       (n_1992), .Q (n_6545));
  AO221X1 g61748(.A (n_5586), .B (n_3223), .C (n_5700), .D (n_3220), .E
       (n_1968), .Q (n_6544));
  AO221X1 g61749(.A (n_5585), .B (n_3223), .C (n_5702), .D (n_3220), .E
       (n_1964), .Q (n_6543));
  AO221X1 g61750(.A (n_5584), .B (n_3223), .C (n_5705), .D (n_3220), .E
       (n_1961), .Q (n_6541));
  AO221X1 g61751(.A (n_5583), .B (n_3223), .C (n_5706), .D (n_3220), .E
       (n_1967), .Q (n_6540));
  NA3X1 g61752(.A (n_3224), .B (n_1977), .C (n_1916), .Q (n_3227));
  AND3X1 g61753(.A (n_3224), .B (n_6238), .C (n_1976), .Q (n_6520));
  AND4X1 g61754(.A (n_3224), .B (n_1977), .C (n_1915), .D (n_5542), .Q
       (n_3226));
  ON21X1 g61755(.A (n_2590), .B (n_1664), .C (n_3224), .Q (n_1662));
  AN21X1 g61756(.A (n_3221), .B (program_counter[1]), .C (n_6218), .Q
       (n_3225));
  NO3X1 g61757(.A (n_6218), .B (n_6595), .C (n_3167), .Q (n_3224));
  NO2X1 g61758(.A (n_3221), .B (n_204), .Q (n_6218));
  INX1 g61759(.A (n_3223), .Q (n_3222));
  NO2X1 g61760(.A (n_3220), .B (n_1848), .Q (n_3223));
  AN21X1 g61762(.A (n_3219), .B (branch_type), .C (n_1806), .Q
       (n_3221));
  NA2X1 g61763(.A (n_3218), .B (n_3216), .Q (n_3219));
  AN21X1 g61764(.A (n_3215), .B (n_6457), .C (n_3217), .Q (n_3218));
  ON211X1 g61765(.A (n_3213), .B (n_1771), .C (n_3214), .D (n_3211), .Q
       (n_3217));
  NA2I1X1 g61766(.B (n_6456), .AN (n_3215), .Q (n_3216));
  ON21X1 g61767(.A (n_3213), .B (n_3114), .C (n_3120), .Q (n_3215));
  NA2X1 g61768(.A (n_3213), .B (n_6454), .Q (n_3214));
  NA2X1 g61769(.A (n_3212), .B (n_1660), .Q (n_3213));
  NA3X1 g61770(.A (n_3210), .B (n_3199), .C (n_3189), .Q (n_3212));
  MU2IX1 g61771(.S (n_3209), .IN0 (n_6459), .IN1 (n_6458), .Q (n_3211));
  ON21X1 g61772(.A (n_3208), .B (n_3192), .C (n_3205), .Q (n_3210));
  NA2X1 g61774(.A (n_1659), .B (n_3204), .Q (n_3209));
  AN21X1 g61775(.A (n_3191), .B (n_3202), .C (n_3201), .Q (n_3208));
  AN22X1 g61777(.A (n_3195), .B (n_3171), .C (n_3194), .D (n_3113), .Q
       (n_3207));
  AN21X1 g61778(.A (n_3196), .B (n_3189), .C (n_3198), .Q (n_3206));
  AN21X1 g61779(.A (n_3197), .B (n_3123), .C (n_3203), .Q (n_3205));
  AND5X1 g61780(.A (n_3200), .B (n_3187), .C (n_3172), .D (n_3154), .E
       (n_3152), .Q (n_3204));
  AN211X1 g61781(.A (n_3186), .B (n_3152), .C (n_3128), .D (n_3175), .Q
       (n_3203));
  ON221X1 g61782(.A (n_3140), .B (n_3184), .C (n_191), .D (n_3092), .E
       (n_3157), .Q (n_3202));
  ON221X1 g61783(.A (n_3094), .B (n_3176), .C (n_3118), .D (n_3153), .E
       (n_3162), .Q (n_3201));
  NO2X1 g61784(.A (n_3192), .B (n_3188), .Q (n_3200));
  NO3X1 g61785(.A (n_3190), .B (n_3173), .C (n_3093), .Q (n_3199));
  ON222X1 g61786(.A (n_3126), .B (n_3148), .C (n_3131), .D (n_3174), .E
       (n_3155), .F (n_3127), .Q (n_3198));
  ON21X1 g61787(.A (n_1656), .B (n_3130), .C (n_3150), .Q (n_3197));
  ON22X1 g61788(.A (n_3146), .B (n_1657), .C (n_3154), .D (n_3124), .Q
       (n_3196));
  ON32X1 g61789(.A (n_3116), .B (n_3151), .C (n_3147), .D (n_3125), .E
       (n_1655), .Q (n_3195));
  ON21X1 g61790(.A (n_1658), .B (n_3097), .C (n_3145), .Q (n_3194));
  AND6X1 g61791(.A (n_3150), .B (n_3126), .C (n_3131), .D (n_3160), .E
       (n_3121), .F (n_3100), .Q (n_3193));
  EO2X1 g61800(.A (alu_2nd_operand[27]), .B (n_1592), .Q (n_6567));
  NA3X1 g61801(.A (n_3168), .B (n_3151), .C (n_3153), .Q (n_3188));
  EO2X1 g61802(.A (alu_2nd_operand[25]), .B (n_1592), .Q (n_6569));
  NO2X1 g61803(.A (n_3173), .B (n_3161), .Q (n_3187));
  EO2X1 g61804(.A (alu_2nd_operand[24]), .B (n_1592), .Q (n_6570));
  AO211X1 g61805(.A (n_3091), .B (n_200), .C (n_3119), .D (n_3156), .Q
       (n_3186));
  EO2X1 g61806(.A (alu_2nd_operand[21]), .B (n_1592), .Q (n_6573));
  EO2X1 g61807(.A (alu_2nd_operand[26]), .B (n_1592), .Q (n_6568));
  EO2X1 g61808(.A (alu_2nd_operand[11]), .B (n_1592), .Q (n_6583));
  EO2X1 g61809(.A (alu_2nd_operand[18]), .B (n_1592), .Q (n_6576));
  EO2X1 g61810(.A (alu_2nd_operand[19]), .B (n_1592), .Q (n_6575));
  EO2X1 g61811(.A (alu_2nd_operand[20]), .B (n_1592), .Q (n_6574));
  OR4X1 g61812(.A (n_3175), .B (n_3144), .C (n_3128), .D (n_3119), .Q
       (n_3192));
  NO2X1 g61813(.A (n_3176), .B (n_3088), .Q (n_3191));
  NA2X1 g61814(.A (n_3171), .B (n_3172), .Q (n_3190));
  NO2X1 g61815(.A (n_3174), .B (n_3102), .Q (n_3189));
  EO2X1 g61816(.A (alu_2nd_operand[16]), .B (n_1592), .Q (n_6578));
  EO2X1 g61817(.A (alu_2nd_operand[10]), .B (n_1592), .Q (n_6584));
  EO2X1 g61818(.A (alu_2nd_operand[23]), .B (n_1592), .Q (n_6571));
  EO2X1 g61819(.A (alu_2nd_operand[22]), .B (n_1592), .Q (n_6572));
  EO2X1 g61820(.A (alu_2nd_operand[14]), .B (n_1592), .Q (n_6580));
  EO2X1 g61821(.A (alu_2nd_operand[15]), .B (n_1592), .Q (n_6579));
  EO2X1 g61822(.A (alu_2nd_operand[28]), .B (n_1592), .Q (n_6566));
  EO2X1 g61823(.A (alu_2nd_operand[30]), .B (n_1592), .Q (n_6564));
  EO2X1 g61824(.A (alu_2nd_operand[6]), .B (n_1592), .Q (n_6588));
  EO2X1 g61826(.A (alu_2nd_operand[29]), .B (n_1592), .Q (n_6565));
  EO2X1 g61827(.A (alu_2nd_operand[31]), .B (n_1592), .Q (n_6563));
  EO2X1 g61828(.A (alu_2nd_operand[9]), .B (n_1592), .Q (n_6585));
  EO2X1 g61829(.A (alu_2nd_operand[12]), .B (n_1592), .Q (n_6582));
  EO2X1 g61830(.A (alu_2nd_operand[8]), .B (n_1592), .Q (n_6586));
  EO2X1 g61831(.A (alu_2nd_operand[13]), .B (n_1592), .Q (n_6581));
  EO2X1 g61832(.A (alu_2nd_operand[17]), .B (n_1592), .Q (n_6577));
  EO2X1 g61833(.A (alu_2nd_operand[7]), .B (n_1592), .Q (n_6587));
  EN2X1 g61834(.A (alu_2nd_operand[5]), .B (n_2076), .Q (n_6589));
  EN2X1 g61835(.A (alu_2nd_operand[4]), .B (n_2076), .Q (n_6590));
  MU2IX1 g61837(.S (n_3139), .IN0 (n_2076), .IN1
       (alu_operation_code_39061), .Q (n_6593));
  AN22X1 g61838(.A (n_3135), .B (n_6729), .C (n_3095), .D (n_6629), .Q
       (n_3184));
  NA2I1X4 g61840(.B (n_3164), .AN (n_3166), .Q (n_6594));
  AN222X1 g61841(.A (n_1907), .B (n_3080), .C (prev_write_data[26]), .D
       (n_1585), .E (n_2263), .F (n_3060), .Q (n_3183));
  AO222X1 g61842(.A (n_3036), .B (n_2382), .C (n_3063), .D (n_2380), .E
       (prev_write_data[14]), .F (n_1585), .Q (write_data[14]));
  AO222X1 g61843(.A (n_3037), .B (n_2382), .C (n_3045), .D (n_2380), .E
       (prev_write_data[13]), .F (n_1585), .Q (write_data[13]));
  AO222X1 g61844(.A (n_3041), .B (n_2382), .C (n_3049), .D (n_2380), .E
       (prev_write_data[12]), .F (n_1585), .Q (write_data[12]));
  AO222X1 g61845(.A (n_3034), .B (n_2382), .C (n_3061), .D (n_2380), .E
       (prev_write_data[11]), .F (n_1585), .Q (write_data[11]));
  AO222X1 g61846(.A (n_3043), .B (n_2382), .C (n_3060), .D (n_2380), .E
       (prev_write_data[10]), .F (n_1585), .Q (write_data[10]));
  AO222X1 g61847(.A (n_3030), .B (n_2382), .C (n_3059), .D (n_2380), .E
       (prev_write_data[9]), .F (n_1585), .Q (write_data[9]));
  AO222X1 g61848(.A (n_3033), .B (n_2382), .C (n_3047), .D (n_2380), .E
       (prev_write_data[8]), .F (n_1585), .Q (write_data[8]));
  AO222X1 g61849(.A (n_1907), .B (n_3076), .C (n_3036), .D (n_2794), .E
       (prev_write_data[22]), .F (n_1585), .Q (write_data[22]));
  AO222X1 g61850(.A (n_1907), .B (n_3056), .C (n_3039), .D (n_2794), .E
       (prev_write_data[23]), .F (n_1585), .Q (write_data[23]));
  AO222X1 g61851(.A (n_1907), .B (n_3082), .C (n_3037), .D (n_2794), .E
       (prev_write_data[21]), .F (n_1585), .Q (write_data[21]));
  AO222X1 g61852(.A (n_1907), .B (n_3085), .C (n_3041), .D (n_2794), .E
       (prev_write_data[20]), .F (n_1585), .Q (write_data[20]));
  AO222X1 g61853(.A (n_1907), .B (n_3065), .C (n_3034), .D (n_2794), .E
       (prev_write_data[19]), .F (n_1585), .Q (write_data[19]));
  AO222X1 g61854(.A (n_1907), .B (n_3054), .C (n_3030), .D (n_2794), .E
       (prev_write_data[17]), .F (n_1585), .Q (write_data[17]));
  AO222X1 g61855(.A (n_1907), .B (n_3057), .C (n_3033), .D (n_2794), .E
       (prev_write_data[16]), .F (n_1585), .Q (write_data[16]));
  AO222X1 g61856(.A (n_1907), .B (n_3068), .C (n_3043), .D (n_2794), .E
       (prev_write_data[18]), .F (n_1585), .Q (write_data[18]));
  AN222X1 g61857(.A (n_1907), .B (n_3084), .C (prev_write_data[31]), .D
       (n_1585), .E (n_2263), .F (n_3062), .Q (n_3182));
  AN222X1 g61858(.A (n_1907), .B (n_3073), .C (prev_write_data[30]), .D
       (n_1585), .E (n_2263), .F (n_3063), .Q (n_3181));
  AN222X1 g61859(.A (n_1907), .B (n_3070), .C (prev_write_data[29]), .D
       (n_1585), .E (n_2263), .F (n_3045), .Q (n_3180));
  AN222X1 g61860(.A (n_1907), .B (n_3072), .C (prev_write_data[28]), .D
       (n_1585), .E (n_2263), .F (n_3049), .Q (n_3179));
  AN222X1 g61861(.A (n_1907), .B (n_3079), .C (prev_write_data[24]), .D
       (n_1585), .E (n_2263), .F (n_3047), .Q (n_3178));
  AN222X1 g61862(.A (n_1907), .B (n_3078), .C (prev_write_data[27]), .D
       (n_1585), .E (n_2263), .F (n_3061), .Q (n_3177));
  AO222X1 g61863(.A (n_3039), .B (n_2382), .C (n_3062), .D (n_2380), .E
       (prev_write_data[15]), .F (n_1585), .Q (write_data[15]));
  AN222X1 g61864(.A (n_1907), .B (n_3067), .C (prev_write_data[25]), .D
       (n_1585), .E (n_2263), .F (n_3059), .Q (n_3170));
  AND3X1 g61865(.A (n_3145), .B (n_3117), .C (n_3115), .Q (n_3169));
  AND2X1 g61866(.A (n_1655), .B (n_3155), .Q (n_3168));
  ON211X1 g61867(.A (n_1990), .B (n_1587), .C (n_2146), .D (n_3132), .Q
       (n_3167));
  NO2X2 g61868(.A (alu_2nd_operand[0]), .B (n_2076), .Q (n_3166));
  NA2X2 g61871(.A (alu_2nd_operand[0]), .B (n_2076), .Q (n_3164));
  NA2X1 g61874(.A (n_3149), .B (n_3098), .Q (n_3162));
  NA3X1 g61876(.A (n_1654), .B (n_3091), .C (n_3094), .Q (n_3161));
  AN211X1 g61877(.A (\rs1_data[0]_39306 ), .B (n_3032), .C (n_3098), .D
       (n_3134), .Q (n_3160));
  NA3I1X1 g61879(.B (n_3096), .C (n_3099), .AN (n_3093), .Q (n_3158));
  AO21X1 g61880(.A (n_3092), .B (n_191), .C (n_3034), .Q (n_3157));
  AN21X1 g61881(.A (n_3090), .B (n_4487), .C (n_1646), .Q (n_3156));
  NA2X1 g61882(.A (n_3149), .B (n_1564), .Q (n_3176));
  NA3I1X1 g61883(.B (n_3143), .C (n_3123), .AN (n_3130), .Q (n_3175));
  OR2X1 g61884(.A (n_3148), .B (n_3110), .Q (n_3174));
  OR2X1 g61885(.A (n_3146), .B (n_3089), .Q (n_3173));
  NO2X1 g61886(.A (n_3147), .B (n_3142), .Q (n_3172));
  NO3X1 g61887(.A (n_3141), .B (n_3097), .C (n_3114), .Q (n_3171));
  AO22X1 g61888(.A (n_2795), .B (n_3039), .C (n_1585), .D
       (prev_write_data[7]), .Q (write_data[7]));
  AO22X1 g61889(.A (n_2795), .B (n_3036), .C (n_1585), .D
       (prev_write_data[6]), .Q (write_data[6]));
  AO22X1 g61890(.A (n_2795), .B (n_3037), .C (n_1585), .D
       (prev_write_data[5]), .Q (write_data[5]));
  AO22X1 g61891(.A (n_2795), .B (n_3041), .C (n_1585), .D
       (prev_write_data[4]), .Q (write_data[4]));
  AO22X1 g61892(.A (n_2795), .B (n_3034), .C (n_1585), .D
       (prev_write_data[3]), .Q (write_data[3]));
  AO22X1 g61893(.A (n_2795), .B (n_3043), .C (n_1585), .D
       (prev_write_data[2]), .Q (write_data[2]));
  AO22X1 g61894(.A (n_2795), .B (n_3030), .C (n_1585), .D
       (prev_write_data[1]), .Q (write_data[1]));
  AO22X1 g61895(.A (n_2795), .B (n_3033), .C (n_1585), .D
       (prev_write_data[0]), .Q (write_data[0]));
  ON22X1 g61896(.A (n_1646), .B (n_4487), .C (\rs1_data[8]_39396 ), .D
       (n_3048), .Q (n_3144));
  NO2X1 g61898(.A (n_3122), .B (n_3103), .Q (n_3143));
  OR2X1 g61899(.A (n_3116), .B (n_3104), .Q (n_3142));
  OR2X1 g61900(.A (n_3129), .B (n_3112), .Q (n_3141));
  AN22X1 g61901(.A (\rs1_data[23]_39246 ), .B (n_3055), .C
       (\rs1_data[22]_39546 ), .D (n_3075), .Q (n_3155));
  AN22X1 g61902(.A (n_3066), .B (n_4477), .C (n_3069), .D (n_4478), .Q
       (n_3154));
  AN22X1 g61903(.A (\rs1_data[7]_39386 ), .B (n_3040), .C (n_4466), .D
       (n_1643), .Q (n_3153));
  AN22X1 g61904(.A (n_1647), .B (n_4480), .C (n_1648), .D (n_4474), .Q
       (n_3152));
  AN22X1 g61905(.A (n_1650), .B (n_4481), .C (n_1651), .D
       (\rs1_data[24]_39256 ), .Q (n_3151));
  AN22X1 g61906(.A (\rs1_data[15]_39476 ), .B (n_1649), .C
       (\rs1_data[14]_39466 ), .D (n_3064), .Q (n_3150));
  NO2X1 g61907(.A (n_3106), .B (n_3118), .Q (n_3149));
  OR2X1 g61909(.A (n_3127), .B (n_3107), .Q (n_3148));
  OR2X1 g61910(.A (n_3111), .B (n_3125), .Q (n_3147));
  OR2X1 g61911(.A (n_3124), .B (n_3109), .Q (n_3146));
  AND2X1 g61912(.A (n_3120), .B (n_3101), .Q (n_3145));
  MU2X1 g61913(.S (\instruction[5]_40139 ), .IN0 (n_6002), .IN1
       (n_3068), .Q (alu_2nd_operand[18]));
  MU2X1 g61914(.S (\instruction[5]_40139 ), .IN0 (n_5992), .IN1
       (n_3085), .Q (alu_2nd_operand[20]));
  MU2X1 g61915(.S (\instruction[5]_40139 ), .IN0 (n_6001), .IN1
       (n_3065), .Q (alu_2nd_operand[19]));
  MU2X1 g61916(.S (\instruction[5]_40139 ), .IN0 (n_5996), .IN1
       (n_3078), .Q (alu_2nd_operand[27]));
  MU2X1 g61917(.S (\instruction[5]_40139 ), .IN0 (n_5997), .IN1
       (n_3080), .Q (alu_2nd_operand[26]));
  MU2X1 g61918(.S (\instruction[5]_40139 ), .IN0 (n_6015), .IN1
       (n_3082), .Q (alu_2nd_operand[21]));
  MU2X1 g61919(.S (\instruction[5]_40139 ), .IN0 (n_6560), .IN1
       (n_3084), .Q (alu_2nd_operand[31]));
  MU2X1 g61920(.S (\instruction[5]_40139 ), .IN0 (n_5993), .IN1
       (n_3073), .Q (alu_2nd_operand[30]));
  MU2X1 g61921(.S (\instruction[5]_40139 ), .IN0 (n_5995), .IN1
       (n_3072), .Q (alu_2nd_operand[28]));
  MU2X1 g61922(.S (\instruction[5]_40139 ), .IN0 (n_5998), .IN1
       (n_3067), .Q (alu_2nd_operand[25]));
  MU2X1 g61923(.S (\instruction[5]_40139 ), .IN0 (n_5999), .IN1
       (n_3079), .Q (alu_2nd_operand[24]));
  MU2X1 g61924(.S (\instruction[5]_40139 ), .IN0 (n_5994), .IN1
       (n_3070), .Q (alu_2nd_operand[29]));
  MU2X1 g61925(.S (\instruction[5]_40139 ), .IN0 (n_6013), .IN1
       (n_3061), .Q (alu_2nd_operand[11]));
  BUX1 g61926(.A (n_3139), .Q (alu_2nd_operand[1]));
  INCX12 g61927(.A (n_3138), .Q (alu_2nd_operand[2]));
  INX8 g61929(.A (n_177), .Q (alu_2nd_operand[3]));
  ON21X1 g61930(.A (n_3051), .B (n_2587), .C (n_121), .Q (n_6486));
  NA3I2X1 g61931(.C (n_3033), .AN (\rs1_data[0]_39306 ), .BN (n_6629),
       .Q (n_3135));
  ON21X1 g61932(.A (n_3059), .B (n_200), .C (n_3095), .Q (n_3134));
  ON21X1 g61933(.A (n_3051), .B (n_2586), .C (n_121), .Q (n_6497));
  ON21X1 g61934(.A (n_3053), .B (n_2589), .C (n_121), .Q (n_6496));
  ON21X1 g61935(.A (n_3052), .B (n_2589), .C (n_121), .Q (n_6495));
  ON21X1 g61936(.A (n_3052), .B (n_2586), .C (n_121), .Q (n_6491));
  ON21X1 g61937(.A (n_3053), .B (n_2586), .C (n_121), .Q (n_6489));
  ON21X1 g61938(.A (n_3051), .B (n_2588), .C (n_121), .Q (n_6488));
  AN22X1 g61939(.A (n_6629), .B (n_6729), .C (n_6757), .D (n_3035), .Q
       (n_3133));
  ON21X1 g61940(.A (n_3052), .B (n_2588), .C (n_121), .Q (n_6484));
  ON21X1 g61941(.A (n_3058), .B (n_2586), .C (n_121), .Q (n_6481));
  ON21X1 g61942(.A (n_3053), .B (n_2588), .C (n_121), .Q (n_6477));
  ON21X1 g61943(.A (n_3052), .B (n_2587), .C (n_121), .Q (n_6475));
  ON21X1 g61944(.A (n_3058), .B (n_2588), .C (n_121), .Q (n_6474));
  ON21X1 g61945(.A (n_3053), .B (n_2587), .C (n_121), .Q (n_6470));
  ON21X1 g61946(.A (n_3051), .B (n_2589), .C (n_121), .Q (n_6468));
  ON21X1 g61947(.A (n_3058), .B (n_2587), .C (n_121), .Q (n_6467));
  OA31X1 g61948(.A (n_1698), .B (n_6453), .C (mret), .D (n_2022), .Q
       (n_3132));
  ON22X1 g61949(.A (n_6628), .B (n_3044), .C (n_6757), .D (n_3035), .Q
       (n_3140));
  MU2IX2 g61950(.S (\instruction[5]_40139 ), .IN0 (n_1702), .IN1
       (n_6729), .Q (n_3139));
  NO2X2 g61951(.A (n_3087), .B (n_1581), .Q (n_3138));
  NA2X4 g61952(.A (n_3086), .B (n_1717), .Q (alu_2nd_operand[0]));
  MU2X1 g61953(.S (\instruction[5]_40139 ), .IN0 (n_6005), .IN1
       (n_3062), .Q (alu_2nd_operand[15]));
  MU2X1 g61954(.S (\instruction[5]_40139 ), .IN0 (n_5991), .IN1
       (n_3076), .Q (alu_2nd_operand[22]));
  MU2X1 g61955(.S (\instruction[5]_40139 ), .IN0 (n_6000), .IN1
       (n_3056), .Q (alu_2nd_operand[23]));
  MU2X1 g61956(.S (\instruction[5]_40139 ), .IN0 (n_6008), .IN1
       (n_3049), .Q (alu_2nd_operand[12]));
  MU2X1 g61957(.S (\instruction[5]_40139 ), .IN0 (n_6557), .IN1
       (n_3047), .Q (alu_2nd_operand[8]));
  OA21X4 g61958(.A (n_3035), .B (n_1686), .C (n_1718), .Q (n_177));
  MU2X1 g61959(.S (\instruction[5]_40139 ), .IN0 (n_6004), .IN1
       (n_3057), .Q (alu_2nd_operand[16]));
  MU2X1 g61960(.S (\instruction[5]_40139 ), .IN0 (n_6555), .IN1
       (n_3036), .Q (alu_2nd_operand[6]));
  MU2X1 g61961(.S (\instruction[5]_40139 ), .IN0 (n_6003), .IN1
       (n_3054), .Q (alu_2nd_operand[17]));
  MU2X1 g61962(.S (\instruction[5]_40139 ), .IN0 (n_6007), .IN1
       (n_3045), .Q (alu_2nd_operand[13]));
  MU2X1 g61963(.S (\instruction[5]_40139 ), .IN0 (n_6559), .IN1
       (n_3060), .Q (alu_2nd_operand[10]));
  MU2X4 g61964(.S (\instruction[5]_40139 ), .IN0 (n_6717), .IN1
       (n_3041), .Q (alu_2nd_operand[4]));
  MU2X1 g61965(.S (\instruction[5]_40139 ), .IN0 (n_6556), .IN1
       (n_3039), .Q (alu_2nd_operand[7]));
  MU2X1 g61966(.S (\instruction[5]_40139 ), .IN0 (n_6554), .IN1
       (n_3037), .Q (alu_2nd_operand[5]));
  MU2X1 g61967(.S (\instruction[5]_40139 ), .IN0 (n_6558), .IN1
       (n_3059), .Q (alu_2nd_operand[9]));
  MU2X1 g61968(.S (\instruction[5]_40139 ), .IN0 (n_6006), .IN1
       (n_3063), .Q (alu_2nd_operand[14]));
  INX1 g61969(.A (n_3114), .Q (n_3113));
  NO2X1 g61970(.A (n_3071), .B (\rs1_data[28]_39296 ), .Q (n_3112));
  NO2X1 g61971(.A (n_3081), .B (\rs1_data[26]_39276 ), .Q (n_3111));
  NO2X1 g61972(.A (n_1652), .B (\rs1_data[21]_39536 ), .Q (n_3110));
  NO2X1 g61973(.A (n_3069), .B (n_4478), .Q (n_3109));
  NA2X1 g61974(.A (\rs1_data[27]_39286 ), .B (n_3077), .Q (n_3108));
  NO2X1 g61975(.A (\rs1_data[22]_39546 ), .B (n_3075), .Q (n_3107));
  NO2X1 g61976(.A (n_4466), .B (n_1643), .Q (n_3106));
  NA2X1 g61977(.A (\rs1_data[26]_39276 ), .B (n_3081), .Q (n_3105));
  NO2X1 g61978(.A (n_1651), .B (\rs1_data[24]_39256 ), .Q (n_3104));
  NO2X1 g61979(.A (n_4475), .B (n_3050), .Q (n_3103));
  NO2I1X1 g61980(.B (n_4486), .AN (n_3085), .Q (n_3102));
  NA2X1 g61981(.A (\rs1_data[30]_39446 ), .B (n_3074), .Q (n_3101));
  NA2X1 g61982(.A (n_1653), .B (n_4486), .Q (n_3131));
  NO2X1 g61983(.A (\rs1_data[14]_39466 ), .B (n_3064), .Q (n_3130));
  NO2I1X1 g61984(.B (\rs1_data[29]_39336 ), .AN (n_3070), .Q (n_3129));
  NO2X1 g61985(.A (n_1648), .B (n_4474), .Q (n_3128));
  NO2X1 g61986(.A (\rs1_data[23]_39246 ), .B (n_3055), .Q (n_3127));
  NA2X1 g61987(.A (n_1652), .B (\rs1_data[21]_39536 ), .Q (n_3126));
  NO2X1 g61988(.A (n_3077), .B (\rs1_data[27]_39286 ), .Q (n_3125));
  NO2X1 g61989(.A (n_3066), .B (n_4477), .Q (n_3124));
  OR2X1 g61990(.A (\rs1_data[15]_39476 ), .B (n_1649), .Q (n_3123));
  NO2X1 g61991(.A (n_4476), .B (n_3046), .Q (n_3122));
  NA2X1 g61992(.A (n_4476), .B (n_3046), .Q (n_3121));
  NA2X1 g61993(.A (n_3083), .B (alu_sra_result[31]), .Q (n_3120));
  NO2X1 g61994(.A (n_1647), .B (n_4480), .Q (n_3119));
  NO2X1 g61995(.A (\rs1_data[7]_39386 ), .B (n_3040), .Q (n_3118));
  NA2I1X1 g61996(.B (\rs1_data[28]_39296 ), .AN (n_3072), .Q (n_3117));
  NO2X1 g61997(.A (n_1650), .B (n_4481), .Q (n_3116));
  NA2I1X1 g61998(.B (\rs1_data[29]_39336 ), .AN (n_3070), .Q (n_3115));
  NO2I1X1 g61999(.B (alu_sra_result[31]), .AN (n_3084), .Q (n_3114));
  INX1 g62000(.A (n_3091), .Q (n_3090));
  AO21X1 g62001(.A (n_2881), .B (n_3024), .C (n_1748), .Q (n_6473));
  NO2X1 g62002(.A (n_1645), .B (\rs1_data[16]_39486 ), .Q (n_3089));
  NO2X1 g62003(.A (n_6627), .B (n_3042), .Q (n_3088));
  ON21X1 g62004(.A (n_2882), .B (n_1576), .C (n_121), .Q (n_6469));
  ON21X1 g62005(.A (n_2886), .B (n_1571), .C (n_121), .Q (n_6471));
  NO2X1 g62007(.A (n_3044), .B (n_1686), .Q (n_3087));
  NA2X4 g62008(.A (n_3033), .B (\instruction[5]_40139 ), .Q (n_3086));
  ON21X1 g62009(.A (n_2886), .B (n_3022), .C (n_121), .Q (n_6498));
  ON21X1 g62010(.A (n_2885), .B (n_3022), .C (n_121), .Q (n_6493));
  AO21X1 g62011(.A (n_2884), .B (n_3024), .C (n_1748), .Q (n_6492));
  ON21X1 g62012(.A (n_2883), .B (n_1571), .C (n_121), .Q (n_6490));
  ON21X1 g62013(.A (n_2886), .B (n_1576), .C (n_121), .Q (n_6494));
  ON21X1 g62014(.A (n_2883), .B (n_3022), .C (n_121), .Q (n_6487));
  ON21X1 g62015(.A (n_2885), .B (n_1576), .C (n_121), .Q (n_6485));
  ON21X1 g62016(.A (n_2882), .B (n_1571), .C (n_121), .Q (n_6483));
  ON21X1 g62017(.A (n_2885), .B (n_1571), .C (n_121), .Q (n_6482));
  ON21X1 g62018(.A (n_2883), .B (n_3023), .C (n_121), .Q (n_6480));
  ON21X1 g62019(.A (n_2882), .B (n_3022), .C (n_121), .Q (n_6478));
  ON21X1 g62020(.A (n_2883), .B (n_1576), .C (n_121), .Q (n_6476));
  ON21X1 g62021(.A (n_2886), .B (n_3023), .C (n_121), .Q (n_6466));
  NA2X1 g62022(.A (n_1645), .B (\rs1_data[16]_39486 ), .Q (n_3100));
  NA2X1 g62023(.A (n_1644), .B (\rs1_data[17]_39496 ), .Q (n_3099));
  AND2X1 g62024(.A (n_3038), .B (n_4461), .Q (n_3098));
  NO2X1 g62025(.A (\rs1_data[30]_39446 ), .B (n_3074), .Q (n_3097));
  NA2X1 g62026(.A (n_4475), .B (n_3050), .Q (n_3096));
  OR2X1 g62027(.A (\rs1_data[0]_39306 ), .B (n_3032), .Q (n_3095));
  NA2X1 g62028(.A (n_6627), .B (n_3042), .Q (n_3094));
  NO2X1 g62029(.A (n_1644), .B (\rs1_data[17]_39496 ), .Q (n_3093));
  NA2X1 g62030(.A (n_6628), .B (n_3044), .Q (n_3092));
  NA2X1 g62031(.A (\rs1_data[8]_39396 ), .B (n_3048), .Q (n_3091));
  INX1 g62032(.A (n_1653), .Q (n_3085));
  INX1 g62033(.A (n_3083), .Q (n_3084));
  INX1 g62034(.A (n_1652), .Q (n_3082));
  INX1 g62035(.A (n_3081), .Q (n_3080));
  INX1 g62036(.A (n_1651), .Q (n_3079));
  INX1 g62037(.A (n_3077), .Q (n_3078));
  INX1 g62038(.A (n_3075), .Q (n_3076));
  INX1 g62039(.A (n_3074), .Q (n_3073));
  INX1 g62040(.A (n_3071), .Q (n_3072));
  INX1 g62041(.A (n_3069), .Q (n_3068));
  INX1 g62042(.A (n_1650), .Q (n_3067));
  INX1 g62043(.A (n_3066), .Q (n_3065));
  INX1 g62044(.A (n_3064), .Q (n_3063));
  INX1 g62045(.A (n_1649), .Q (n_3062));
  INX1 g62046(.A (n_1648), .Q (n_3061));
  INX1 g62047(.A (n_1647), .Q (n_3060));
  INX1 g62048(.A (n_1646), .Q (n_3059));
  AND5X1 g62051(.A (n_1635), .B (n_2938), .C (n_2920), .D (n_2933), .E
       (n_2930), .Q (n_3083));
  NO2X1 g62053(.A (n_3027), .B (n_2998), .Q (n_3081));
  NO2X1 g62055(.A (n_3026), .B (n_3025), .Q (n_3077));
  NO2X1 g62056(.A (n_3021), .B (n_3018), .Q (n_3075));
  AND5X1 g62057(.A (n_1636), .B (n_2932), .C (n_2929), .D (n_2908), .E
       (n_2953), .Q (n_3074));
  NO2X1 g62058(.A (n_3028), .B (n_3019), .Q (n_3071));
  NA2X1 g62059(.A (n_1637), .B (n_1632), .Q (n_3070));
  AND5X1 g62060(.A (n_1628), .B (n_2940), .C (n_2919), .D (n_2918), .E
       (n_2861), .Q (n_3069));
  AND5X1 g62062(.A (n_1626), .B (n_2912), .C (n_2891), .D (n_2902), .E
       (n_2905), .Q (n_3066));
  AND2X1 g62063(.A (n_1639), .B (n_1627), .Q (n_3064));
  INX1 g62068(.A (n_1645), .Q (n_3057));
  INX1 g62069(.A (n_3055), .Q (n_3056));
  INX1 g62070(.A (n_1644), .Q (n_3054));
  INX1 g62071(.A (n_3050), .Q (n_3049));
  INX1 g62072(.A (n_3048), .Q (n_3047));
  INX1 g62073(.A (n_3046), .Q (n_3045));
  INX1 g62074(.A (n_3044), .Q (n_3043));
  INX2 g62075(.A (n_3042), .Q (n_3041));
  INX1 g62076(.A (n_3040), .Q (n_3039));
  INX1 g62077(.A (n_3038), .Q (n_3037));
  INX1 g62078(.A (n_1643), .Q (n_3036));
  INX1 g62079(.A (n_3035), .Q (n_3034));
  INX1 g62080(.A (n_3033), .Q (n_3032));
  INX1 g62081(.A (n_6729), .Q (n_3030));
  AND3X1 g62082(.A (n_5724), .B (n_2996), .C (n_1813), .Q (n_6217));
  NO6I2X1 g62083(.C (n_6596), .D (n_1772), .E (n_1753), .F
       (instruction[26]), .AN (n_1820), .BN (n_1757), .Q (mret));
  OR2X1 g62084(.A (n_2323), .B (n_1576), .Q (n_3058));
  NO2X1 g62086(.A (n_3020), .B (n_3017), .Q (n_3055));
  NA2X1 g62088(.A (n_2322), .B (n_3024), .Q (n_3053));
  OR2X1 g62089(.A (n_2323), .B (n_3022), .Q (n_3052));
  OR2X1 g62090(.A (n_2323), .B (n_1571), .Q (n_3051));
  NO2X1 g62091(.A (n_3012), .B (n_3016), .Q (n_3050));
  NO2X1 g62092(.A (n_3011), .B (n_3015), .Q (n_3048));
  NO2X1 g62093(.A (n_3013), .B (n_3014), .Q (n_3046));
  NO2X4 g62094(.A (n_3000), .B (n_3002), .Q (n_3044));
  NO2X4 g62095(.A (n_3010), .B (n_3008), .Q (n_3042));
  NO2X1 g62096(.A (n_3006), .B (n_3009), .Q (n_3040));
  NO2X4 g62099(.A (n_3007), .B (n_3005), .Q (n_3035));
  NA2X4 g62100(.A (n_2999), .B (n_3001), .Q (n_3033));
  NA2X4 g62103(.A (n_2994), .B (n_1805), .Q (n_5988));
  NA2X4 g62104(.A (n_2992), .B (n_1811), .Q (n_5987));
  AO22X1 g62105(.A (n_1903), .B (csr_data_out[26]), .C
       (\rs1_data[26]_39276 ), .D (n_1586), .Q (n_5733));
  AO22X2 g62106(.A (n_1886), .B (csr_data_out[30]), .C
       (\rs1_data[30]_39446 ), .D (n_1586), .Q (n_5729));
  AO22X2 g62108(.A (n_1897), .B (csr_data_out[31]), .C
       (alu_sra_result[31]), .D (n_1586), .Q (n_5985));
  AO22X2 g62109(.A (n_1896), .B (csr_data_out[29]), .C
       (\rs1_data[29]_39336 ), .D (n_1586), .Q (n_5730));
  AO22X2 g62110(.A (n_1895), .B (csr_data_out[28]), .C
       (\rs1_data[28]_39296 ), .D (n_1586), .Q (n_5731));
  AO22X2 g62111(.A (n_1898), .B (csr_data_out[27]), .C
       (\rs1_data[27]_39286 ), .D (n_1586), .Q (n_5732));
  AO22X1 g62112(.A (n_1893), .B (csr_data_out[23]), .C
       (\rs1_data[23]_39246 ), .D (n_1586), .Q (n_5736));
  AO22X2 g62113(.A (n_1892), .B (csr_data_out[22]), .C
       (\rs1_data[22]_39546 ), .D (n_1586), .Q (n_5737));
  AO22X1 g62114(.A (n_1891), .B (csr_data_out[15]), .C
       (\rs1_data[15]_39476 ), .D (n_1586), .Q (n_4538));
  AO22X1 g62115(.A (n_1894), .B (csr_data_out[14]), .C
       (\rs1_data[14]_39466 ), .D (n_1586), .Q (n_4536));
  AO22X2 g62116(.A (n_1889), .B (csr_data_out[21]), .C
       (\rs1_data[21]_39536 ), .D (n_1586), .Q (n_5738));
  AO22X2 g62117(.A (n_1888), .B (csr_data_out[19]), .C (n_4477), .D
       (n_1586), .Q (n_5740));
  AO22X2 g62118(.A (n_1887), .B (csr_data_out[18]), .C (n_4478), .D
       (n_1586), .Q (n_5741));
  AO22X2 g62119(.A (n_1890), .B (csr_data_out[11]), .C (n_4474), .D
       (n_1586), .Q (n_5748));
  AO22X1 g62120(.A (n_1885), .B (csr_data_out[25]), .C (n_4481), .D
       (n_1586), .Q (n_5734));
  AO22X2 g62121(.A (n_1884), .B (csr_data_out[24]), .C
       (\rs1_data[24]_39256 ), .D (n_1586), .Q (n_5735));
  AO22X2 g62122(.A (n_1881), .B (csr_data_out[20]), .C (n_4486), .D
       (n_1586), .Q (n_5739));
  AO22X2 g62123(.A (n_1883), .B (csr_data_out[13]), .C (n_4476), .D
       (n_1586), .Q (n_5746));
  AO22X2 g62124(.A (n_1882), .B (csr_data_out[12]), .C (n_4475), .D
       (n_1586), .Q (n_5747));
  AO22X1 g62125(.A (n_1880), .B (csr_data_out[10]), .C (n_4480), .D
       (n_1586), .Q (n_5749));
  AO22X1 g62127(.A (n_1875), .B (csr_data_out[16]), .C
       (\rs1_data[16]_39486 ), .D (n_1586), .Q (n_5743));
  AO22X2 g62128(.A (n_1876), .B (csr_data_out[8]), .C
       (\rs1_data[8]_39396 ), .D (n_1586), .Q (n_5751));
  AO22X1 g62129(.A (n_1874), .B (csr_data_out[9]), .C (n_4487), .D
       (n_1586), .Q (n_5750));
  AO22X2 g62131(.A (n_1872), .B (csr_data_out[17]), .C
       (\rs1_data[17]_39496 ), .D (n_1586), .Q (n_5742));
  NA3X1 g62132(.A (n_2989), .B (n_2941), .C (n_2923), .Q (n_3028));
  NA3X1 g62133(.A (n_2990), .B (n_2939), .C (n_2915), .Q (n_3027));
  NA3X1 g62135(.A (n_2988), .B (n_2937), .C (n_2921), .Q (n_3026));
  NA3X1 g62138(.A (n_2995), .B (n_1617), .C (n_1618), .Q (n_3025));
  AO22X2 g62143(.A (n_1904), .B (csr_data_out[4]), .C (n_1775), .D
       (n_1767), .Q (n_4535));
  INX1 g62144(.A (n_3024), .Q (n_3023));
  NA3X1 g62145(.A (n_2985), .B (n_2897), .C (n_2901), .Q (n_3021));
  NA3X1 g62146(.A (n_2984), .B (n_2900), .C (n_2896), .Q (n_3020));
  NA3X1 g62153(.A (n_2982), .B (n_2904), .C (n_2903), .Q (n_3019));
  NA3X1 g62157(.A (n_2981), .B (n_1620), .C (n_2845), .Q (n_3018));
  NA3X1 g62158(.A (n_2980), .B (n_2946), .C (n_2844), .Q (n_3017));
  NA3X1 g62159(.A (n_2975), .B (n_6734), .C (n_6748), .Q (n_3016));
  NA3X1 g62160(.A (n_2974), .B (n_1613), .C (n_1612), .Q (n_3015));
  NA3X1 g62161(.A (n_2976), .B (n_6736), .C (n_6735), .Q (n_3014));
  NA3X1 g62163(.A (n_2986), .B (n_2895), .C (n_2851), .Q (n_3013));
  NA3X1 g62164(.A (n_2969), .B (n_2931), .C (n_2850), .Q (n_3012));
  NA3X1 g62165(.A (n_2977), .B (n_1619), .C (n_6744), .Q (n_3011));
  NA3X1 g62167(.A (n_2973), .B (n_2824), .C (n_2823), .Q (n_3010));
  NA3X1 g62169(.A (n_2970), .B (n_2854), .C (n_1611), .Q (n_3009));
  NA3X1 g62171(.A (n_2967), .B (n_1608), .C (n_2807), .Q (n_3008));
  NA2X1 g62172(.A (n_2978), .B (n_2972), .Q (n_3007));
  NA3X1 g62174(.A (n_2971), .B (n_2847), .C (n_2857), .Q (n_3006));
  NA3X2 g62175(.A (n_6760), .B (n_2833), .C (n_2834), .Q (n_3005));
  NA3X1 g62177(.A (n_2965), .B (n_6752), .C (n_6755), .Q (n_3003));
  NA3X1 g62178(.A (n_2961), .B (n_2799), .C (n_2808), .Q (n_3002));
  NO3X2 g62179(.A (n_6733), .B (n_2798), .C (n_2818), .Q (n_3001));
  NA3X1 g62180(.A (n_2962), .B (n_1605), .C (n_1604), .Q (n_3000));
  NO3X4 g62181(.A (n_2963), .B (n_2805), .C (n_2803), .Q (n_2999));
  NA3X1 g62182(.A (n_2987), .B (n_6738), .C (n_2860), .Q (n_2998));
  NO2X1 g62183(.A (n_2997), .B (n_1769), .Q (n_3024));
  NA2X1 g62185(.A (n_2997), .B (n_1769), .Q (n_3022));
  INX1 g62188(.A (n_2996), .Q (n_6596));
  HAX1 g62189(.A (n_2379), .B (n_1701), .S (n_2997), .CO (n_2996));
  NO2X1 g62190(.A (n_2909), .B (n_2952), .Q (n_2995));
  NA2X1 g62191(.A (n_1861), .B (csr_data_out[2]), .Q (n_2994));
  NA2X1 g62193(.A (n_1900), .B (csr_data_out[3]), .Q (n_2992));
  AND4X1 g62195(.A (n_2737), .B (n_2744), .C (n_2736), .D (n_2749), .Q
       (n_2990));
  NO2X1 g62196(.A (n_2907), .B (n_6737), .Q (n_2989));
  NO2X1 g62197(.A (n_2922), .B (n_6743), .Q (n_2988));
  AND4X1 g62198(.A (n_2667), .B (n_2669), .C (n_2668), .D (n_2521), .Q
       (n_2987));
  NO2X1 g62199(.A (n_6785), .B (n_6740), .Q (n_2986));
  AND4X1 g62200(.A (n_2635), .B (n_2677), .C (n_2692), .D (n_2694), .Q
       (n_2985));
  AND4X1 g62201(.A (n_2631), .B (n_2673), .C (n_2793), .D (n_2693), .Q
       (n_2984));
  AND3X1 g62202(.A (n_6745), .B (n_2700), .C (n_2617), .Q (n_2983));
  AND4X1 g62203(.A (n_2600), .B (n_2599), .C (n_2601), .D (n_2499), .Q
       (n_2982));
  AND4X1 g62204(.A (n_2591), .B (n_2593), .C (n_2592), .D (n_2480), .Q
       (n_2981));
  AND4X1 g62205(.A (n_2584), .B (n_2791), .C (n_2482), .D (n_2479), .Q
       (n_2980));
  AND4X1 g62206(.A (n_2583), .B (n_2581), .C (n_2582), .D (n_2478), .Q
       (n_2979));
  OR2X1 g62207(.A (n_6215), .B (n_6216), .Q (n_6595));
  NO2X1 g62208(.A (n_2816), .B (n_2806), .Q (n_2978));
  NO2X1 g62209(.A (n_2875), .B (n_2830), .Q (n_2977));
  NO2X1 g62210(.A (n_2836), .B (n_6750), .Q (n_2976));
  AND4X1 g62211(.A (n_2506), .B (n_2508), .C (n_2507), .D (n_2462), .Q
       (n_2975));
  AND4X1 g62212(.A (n_2500), .B (n_2502), .C (n_2501), .D (n_2461), .Q
       (n_2974));
  AND4X1 g62213(.A (n_2465), .B (n_2467), .C (n_2466), .D (n_2468), .Q
       (n_2973));
  NO2X1 g62214(.A (n_2838), .B (n_2815), .Q (n_2972));
  NO2X1 g62215(.A (n_2852), .B (n_2813), .Q (n_2971));
  AND4X1 g62216(.A (n_2452), .B (n_2454), .C (n_2453), .D (n_2421), .Q
       (n_2970));
  NO2X1 g62217(.A (n_6741), .B (n_6749), .Q (n_2969));
  AND4X1 g62219(.A (n_2439), .B (n_2441), .C (n_2440), .D (n_2417), .Q
       (n_2967));
  NO2X1 g62221(.A (n_2802), .B (n_2800), .Q (n_2965));
  NA3X2 g62223(.A (n_6754), .B (n_2410), .C (n_2388), .Q (n_2963));
  NO2X1 g62224(.A (n_2804), .B (n_6747), .Q (n_2962));
  AND4X1 g62225(.A (n_2393), .B (n_2398), .C (n_2394), .D (n_2386), .Q
       (n_2961));
  NA6X1 g62226(.A (n_2304), .B (n_2039), .C (n_2034), .D (n_2040), .E
       (n_2131), .F (n_2130), .Q (csr_data_out[7]));
  OR2X1 g62228(.A (n_2794), .B (n_1907), .Q (n_2959));
  AND2X1 g62231(.A (n_2579), .B (n_2580), .Q (n_2956));
  AN222X1 g62232(.A (n_2159), .B (n_4592), .C (n_4584), .D (n_1595), .E
       (n_4581), .F (n_2188), .Q (n_2955));
  AN221X1 g62234(.A (n_5199), .B (n_2173), .C (n_5198), .D (n_1600), .E
       (n_2520), .Q (n_2953));
  NA2X1 g62235(.A (n_2672), .B (n_2522), .Q (n_2952));
  AN221X1 g62236(.A (n_5540), .B (n_2173), .C (n_5539), .D (n_1600), .E
       (n_2523), .Q (n_2951));
  AN221X1 g62237(.A (n_5474), .B (n_2171), .C (n_5473), .D (n_2167), .E
       (n_2524), .Q (n_2950));
  AN221X1 g62238(.A (n_5137), .B (n_2173), .C (n_5132), .D (n_2167), .E
       (n_2525), .Q (n_2949));
  AN221X1 g62239(.A (n_5443), .B (n_2171), .C (n_5442), .D (n_2167), .E
       (n_2543), .Q (n_2948));
  AN221X1 g62240(.A (n_5420), .B (n_2185), .C (n_5419), .D (n_2187), .E
       (n_2765), .Q (n_2947));
  AND2X1 g62241(.A (n_2625), .B (n_2675), .Q (n_2946));
  AN222X1 g62243(.A (n_2159), .B (n_5429), .C (n_5425), .D (n_2160), .E
       (n_5430), .F (n_2164), .Q (n_2945));
  AN221X1 g62244(.A (n_5296), .B (n_2185), .C (n_5295), .D (n_2187), .E
       (n_2574), .Q (n_2944));
  AN221X1 g62245(.A (n_5327), .B (n_2185), .C (n_5326), .D (n_2187), .E
       (n_2575), .Q (n_2943));
  AN221X1 g62247(.A (n_5451), .B (n_2185), .C (n_5450), .D (n_2187), .E
       (n_2773), .Q (n_2942));
  AND2X1 g62248(.A (n_2782), .B (n_2772), .Q (n_2941));
  AN221X1 g62249(.A (n_5358), .B (n_2185), .C (n_5357), .D (n_2187), .E
       (n_2769), .Q (n_2940));
  AND2X1 g62250(.A (n_2780), .B (n_2768), .Q (n_2939));
  AN221X1 g62251(.A (n_5517), .B (n_2200), .C (n_5519), .D (n_2153), .E
       (n_2771), .Q (n_2938));
  AND2X1 g62252(.A (n_2762), .B (n_2770), .Q (n_2937));
  AN221X1 g62253(.A (n_5424), .B (n_2200), .C (n_5426), .D (n_2153), .E
       (n_2754), .Q (n_2936));
  AN221X1 g62254(.A (n_5435), .B (n_2179), .C (n_5434), .D (n_2177), .E
       (n_2757), .Q (n_2935));
  AN221X1 g62255(.A (n_5471), .B (n_2191), .C (n_5467), .D (n_2183), .E
       (n_2752), .Q (n_2934));
  AN221X1 g62256(.A (n_5533), .B (n_2191), .C (n_5529), .D (n_2183), .E
       (n_2740), .Q (n_2933));
  AN221X1 g62258(.A (n_5192), .B (n_2191), .C (n_5188), .D (n_2183), .E
       (n_2748), .Q (n_2932));
  AND2X1 g62259(.A (n_2577), .B (n_2570), .Q (n_2931));
  AN221X1 g62261(.A (n_5526), .B (n_2181), .C (n_5528), .D (n_2179), .E
       (n_2750), .Q (n_2930));
  AN221X1 g62262(.A (n_5185), .B (n_2181), .C (n_5186), .D (n_2177), .E
       (n_2735), .Q (n_2929));
  AN221X1 g62263(.A (n_4586), .B (n_2202), .C (n_4585), .D (n_2198), .E
       (n_2734), .Q (n_2928));
  AND2X1 g62264(.A (n_2777), .B (n_2733), .Q (n_2927));
  AN221X1 g62265(.A (n_5111), .B (n_1596), .C (n_5108), .D (n_2188), .E
       (n_2731), .Q (n_2926));
  AN221X1 g62266(.A (n_5114), .B (n_2200), .C (n_5116), .D (n_2153), .E
       (n_2730), .Q (n_2925));
  AN221X1 g62267(.A (n_5455), .B (n_2200), .C (n_5457), .D (n_2153), .E
       (n_2727), .Q (n_2924));
  AN221X1 g62268(.A (n_4711), .B (n_2200), .C (n_4713), .D (n_2153), .E
       (n_2725), .Q (n_2923));
  NA2X1 g62269(.A (n_2788), .B (n_2723), .Q (n_2922));
  AND2X1 g62270(.A (n_2781), .B (n_2722), .Q (n_2921));
  AN221X1 g62271(.A (n_5513), .B (n_2185), .C (n_5512), .D (n_2187), .E
       (n_2713), .Q (n_2920));
  AN221X1 g62272(.A (n_5359), .B (n_1595), .C (n_5356), .D (n_2188), .E
       (n_2721), .Q (n_2919));
  AN221X1 g62273(.A (n_5362), .B (n_2200), .C (n_5364), .D (n_2153), .E
       (n_2720), .Q (n_2918));
  AND2X1 g62276(.A (n_2761), .B (n_2717), .Q (n_2915));
  AN221X1 g62277(.A (n_4615), .B (n_1596), .C (n_4612), .D (n_2188), .E
       (n_2716), .Q (n_2914));
  AN221X1 g62278(.A (n_4617), .B (n_2202), .C (n_4616), .D (n_2198), .E
       (n_2714), .Q (n_2913));
  AN221X1 g62279(.A (n_5389), .B (n_2185), .C (n_5388), .D (n_2187), .E
       (n_2701), .Q (n_2912));
  AN221X1 g62280(.A (n_5265), .B (n_2185), .C (n_5264), .D (n_2187), .E
       (n_2699), .Q (n_2911));
  AND2X1 g62281(.A (n_2681), .B (n_2682), .Q (n_2910));
  NA2X1 g62282(.A (n_2670), .B (n_2671), .Q (n_2909));
  AN221X1 g62283(.A (n_5197), .B (n_2165), .C (n_5194), .D (n_2167), .E
       (n_2666), .Q (n_2908));
  NA2X1 g62284(.A (n_2726), .B (n_2612), .Q (n_2907));
  AN221X1 g62285(.A (n_4595), .B (n_2154), .C (n_4588), .D (n_2160), .E
       (n_2611), .Q (n_2906));
  AN221X1 g62286(.A (n_5406), .B (n_2193), .C (n_5407), .D (n_2195), .E
       (n_2650), .Q (n_2905));
  AND2X1 g62287(.A (n_2686), .B (n_2653), .Q (n_2904));
  AN221X1 g62288(.A (n_4720), .B (n_2181), .C (n_4725), .D (n_2195), .E
       (n_2652), .Q (n_2903));
  AN221X1 g62289(.A (n_5404), .B (n_2179), .C (n_5403), .D (n_2177), .E
       (n_2651), .Q (n_2902));
  AND2X1 g62290(.A (n_2642), .B (n_2632), .Q (n_2901));
  AND2X1 g62291(.A (n_2641), .B (n_2630), .Q (n_2900));
  AND2X1 g62292(.A (n_2640), .B (n_2627), .Q (n_2899));
  AND2X1 g62293(.A (n_2639), .B (n_2626), .Q (n_2898));
  AND2X1 g62294(.A (n_2634), .B (n_2633), .Q (n_2897));
  AND2X1 g62295(.A (n_2629), .B (n_2628), .Q (n_2896));
  AND2X1 g62296(.A (n_2578), .B (n_2572), .Q (n_2895));
  AND2X1 g62297(.A (n_2594), .B (n_2595), .Q (n_2894));
  AND2X1 g62298(.A (n_2597), .B (n_2598), .Q (n_2893));
  AND2X1 g62300(.A (n_2705), .B (n_2623), .Q (n_2892));
  AN221X1 g62302(.A (n_5393), .B (n_2200), .C (n_5395), .D (n_2153), .E
       (n_2619), .Q (n_2891));
  AND2X1 g62303(.A (n_2698), .B (n_2616), .Q (n_2890));
  AND2X1 g62305(.A (n_2608), .B (n_2610), .Q (n_2889));
  AN221X1 g62306(.A (n_4856), .B (n_2165), .C (n_4857), .D (n_1600), .E
       (n_2607), .Q (n_2888));
  AND2X1 g62307(.A (n_2605), .B (n_2606), .Q (n_2887));
  NA6X1 g62308(.A (n_2141), .B (n_2142), .C (n_2050), .D (n_2049), .E
       (n_2008), .F (n_2037), .Q (csr_data_out[12]));
  NA6X1 g62309(.A (n_2252), .B (n_2139), .C (n_2138), .D (n_2007), .E
       (n_2136), .F (n_2035), .Q (csr_data_out[11]));
  NA3X1 g62310(.A (n_2251), .B (n_2371), .C (n_2047), .Q
       (csr_data_out[10]));
  NA3X1 g62311(.A (n_2254), .B (n_2374), .C (n_2051), .Q
       (csr_data_out[13]));
  NA3X1 g62312(.A (n_2253), .B (n_2373), .C (n_2054), .Q
       (csr_data_out[14]));
  NA3X1 g62313(.A (n_2255), .B (n_2375), .C (n_2055), .Q
       (csr_data_out[15]));
  NA6X1 g62314(.A (n_2101), .B (n_2215), .C (n_2061), .D (n_2072), .E
       (n_2261), .F (n_2143), .Q (csr_data_out[16]));
  NA6X1 g62315(.A (n_2097), .B (n_2232), .C (n_2058), .D (n_2073), .E
       (n_2216), .F (n_2144), .Q (csr_data_out[17]));
  NA6X1 g62316(.A (n_2098), .B (n_2233), .C (n_2062), .D (n_2074), .E
       (n_2218), .F (n_2145), .Q (csr_data_out[18]));
  NA6X1 g62317(.A (n_2099), .B (n_2234), .C (n_2063), .D (n_2105), .E
       (n_2219), .F (n_2259), .Q (csr_data_out[19]));
  NA6X1 g62318(.A (n_2100), .B (n_2244), .C (n_2057), .D (n_2043), .E
       (n_2217), .F (n_2120), .Q (csr_data_out[20]));
  NA6X1 g62319(.A (n_2096), .B (n_2235), .C (n_2059), .D (n_2116), .E
       (n_2220), .F (n_2260), .Q (csr_data_out[21]));
  NA6X1 g62320(.A (n_2095), .B (n_2238), .C (n_2067), .D (n_2112), .E
       (n_2224), .F (n_2258), .Q (csr_data_out[25]));
  NA6X1 g62321(.A (n_2094), .B (n_2246), .C (n_2064), .D (n_2115), .E
       (n_2221), .F (n_2257), .Q (csr_data_out[22]));
  NA6X1 g62322(.A (n_2090), .B (n_2236), .C (n_2065), .D (n_2114), .E
       (n_2222), .F (n_2231), .Q (csr_data_out[23]));
  NA6X1 g62323(.A (n_2093), .B (n_2237), .C (n_2066), .D (n_2113), .E
       (n_2223), .F (n_2206), .Q (csr_data_out[24]));
  NA6X1 g62324(.A (n_2092), .B (n_2239), .C (n_2070), .D (n_2111), .E
       (n_2225), .F (n_2207), .Q (csr_data_out[26]));
  NA6X1 g62325(.A (n_2088), .B (n_2240), .C (n_2068), .D (n_2110), .E
       (n_2226), .F (n_2210), .Q (csr_data_out[27]));
  NA6X1 g62326(.A (n_2087), .B (n_2241), .C (n_2060), .D (n_2109), .E
       (n_2229), .F (n_2211), .Q (csr_data_out[28]));
  NA6X1 g62327(.A (n_2089), .B (n_2242), .C (n_2069), .D (n_2108), .E
       (n_2227), .F (n_2212), .Q (csr_data_out[29]));
  NA6X1 g62328(.A (n_2256), .B (n_2243), .C (n_1997), .D (n_2247), .E
       (n_2213), .F (n_2046), .Q (csr_data_out[30]));
  NA6X1 g62329(.A (n_2091), .B (n_2245), .C (n_2071), .D (n_2106), .E
       (n_2228), .F (n_2214), .Q (csr_data_out[31]));
  NO3X1 g62330(.A (n_2796), .B (n_1948), .C (n_6367), .Q (n_6216));
  AND3X1 g62331(.A (n_2797), .B (n_1768), .C (store_type), .Q (n_6215));
  INX1 g62332(.A (n_2884), .Q (n_2885));
  INX1 g62333(.A (n_2881), .Q (n_2882));
  AN221X1 g62337(.A (n_5315), .B (n_2196), .C (n_5314), .D (n_2195), .E
       (n_2550), .Q (n_2879));
  AN221X1 g62338(.A (n_5309), .B (n_2181), .C (n_5310), .D (n_2177), .E
       (n_2549), .Q (n_2878));
  NA2X1 g62341(.A (n_2569), .B (n_2535), .Q (n_2875));
  AN221X1 g62342(.A (n_5328), .B (n_1596), .C (n_5325), .D (n_2188), .E
       (n_2533), .Q (n_2874));
  AN221X1 g62343(.A (n_4604), .B (n_2169), .C (n_4605), .D (n_2167), .E
       (n_2512), .Q (n_2873));
  AN221X1 g62344(.A (n_4854), .B (n_2171), .C (n_4853), .D (n_2167), .E
       (n_2505), .Q (n_2872));
  AN221X1 g62345(.A (n_5106), .B (n_2173), .C (n_5105), .D (n_1600), .E
       (n_2504), .Q (n_2871));
  AN221X1 g62347(.A (n_5381), .B (n_2171), .C (n_5380), .D (n_2167), .E
       (n_2497), .Q (n_2869));
  AN221X1 g62348(.A (n_4635), .B (n_2169), .C (n_4636), .D (n_2167), .E
       (n_2493), .Q (n_2868));
  AN221X1 g62349(.A (n_5416), .B (n_2173), .C (n_5415), .D (n_1598), .E
       (n_2498), .Q (n_2867));
  AN222X1 g62350(.A (n_2159), .B (n_4840), .C (n_4836), .D (n_2160), .E
       (n_4841), .F (n_2164), .Q (n_2866));
  AN221X1 g62351(.A (n_5518), .B (n_2160), .C (n_5523), .D (n_2164), .E
       (n_2369), .Q (n_2865));
  AN222X1 g62352(.A (n_2159), .B (n_5119), .C (n_5115), .D (n_2160), .E
       (n_5120), .F (n_2164), .Q (n_2864));
  AN221X1 g62353(.A (n_5456), .B (n_2160), .C (n_5461), .D (n_2164), .E
       (n_2368), .Q (n_2863));
  AN222X1 g62355(.A (n_2159), .B (n_5367), .C (n_5363), .D (n_2160), .E
       (n_5368), .F (n_2164), .Q (n_2861));
  AN222X1 g62356(.A (n_2159), .B (n_4654), .C (n_4650), .D (n_2160), .E
       (n_4655), .F (n_2164), .Q (n_2860));
  AN221X1 g62357(.A (n_5177), .B (n_2160), .C (n_5182), .D (n_2164), .E
       (n_2366), .Q (n_2859));
  AN222X1 g62358(.A (n_2159), .B (n_4623), .C (n_4619), .D (n_2160), .E
       (n_4624), .F (n_2164), .Q (n_2858));
  AND2X1 g62359(.A (n_2481), .B (n_2472), .Q (n_2857));
  AN221X1 g62360(.A (n_4939), .B (n_2179), .C (n_4938), .D (n_2177), .E
       (n_2489), .Q (n_2856));
  AN221X1 g62361(.A (n_4943), .B (n_2196), .C (n_4937), .D (n_2181), .E
       (n_2488), .Q (n_2855));
  AND2X1 g62362(.A (n_2483), .B (n_2491), .Q (n_2854));
  AN221X1 g62364(.A (n_5057), .B (n_2159), .C (n_5046), .D (n_2188), .E
       (n_2365), .Q (n_2853));
  NA2X1 g62365(.A (n_2514), .B (n_2473), .Q (n_2852));
  NA2X1 g62366(.A (n_2590), .B (n_1585), .Q (n_6463));
  AND2X1 g62367(.A (n_2548), .B (n_2540), .Q (n_2851));
  AND2X1 g62368(.A (n_2547), .B (n_2537), .Q (n_2850));
  AN221X1 g62370(.A (n_4924), .B (n_2185), .C (n_4923), .D (n_2187), .E
       (n_2515), .Q (n_2848));
  AND2X1 g62371(.A (n_2513), .B (n_2517), .Q (n_2847));
  AN221X1 g62372(.A (n_5259), .B (n_2165), .C (n_5260), .D (n_1600), .E
       (n_2477), .Q (n_2846));
  AN221X1 g62373(.A (n_5487), .B (n_2160), .C (n_5492), .D (n_2164), .E
       (n_2358), .Q (n_2845));
  AN221X1 g62374(.A (n_4557), .B (n_2160), .C (n_4562), .D (n_2164), .E
       (n_2357), .Q (n_2844));
  AN222X1 g62375(.A (n_2159), .B (n_5088), .C (n_5084), .D (n_2160), .E
       (n_5089), .F (n_2164), .Q (n_2843));
  AN221X1 g62376(.A (n_5394), .B (n_2160), .C (n_5399), .D (n_2164), .E
       (n_2363), .Q (n_2842));
  AN221X1 g62378(.A (n_5239), .B (n_2160), .C (n_5244), .D (n_2164), .E
       (n_2360), .Q (n_2840));
  NA2X1 g62381(.A (n_2449), .B (n_2448), .Q (n_2838));
  NA2X1 g62383(.A (n_2509), .B (n_2510), .Q (n_2836));
  AN221X1 g62384(.A (n_5352), .B (n_2165), .C (n_5354), .D (n_2173), .E
       (n_2496), .Q (n_2835));
  NO2X1 g62385(.A (n_2443), .B (n_2444), .Q (n_2834));
  NA2X1 g62389(.A (n_2536), .B (n_2349), .Q (n_2830));
  AN222X1 g62390(.A (n_2159), .B (n_5336), .C (n_5332), .D (n_2160), .E
       (n_5337), .F (n_2164), .Q (n_2829));
  AN221X1 g62391(.A (n_5301), .B (n_2160), .C (n_5306), .D (n_2164), .E
       (n_2343), .Q (n_2828));
  AN221X1 g62394(.A (n_5350), .B (n_2171), .C (n_5349), .D (n_2167), .E
       (n_2460), .Q (n_2826));
  AN221X1 g62395(.A (n_5323), .B (n_2173), .C (n_5322), .D (n_1598), .E
       (n_2459), .Q (n_2825));
  AND2X1 g62397(.A (n_2469), .B (n_2463), .Q (n_2824));
  AN221X1 g62398(.A (n_4901), .B (n_2150), .C (n_4900), .D (n_2152), .E
       (n_2471), .Q (n_2823));
  AND2X1 g62401(.A (n_2455), .B (n_2456), .Q (n_2821));
  NA2X1 g62402(.A (n_2429), .B (n_2430), .Q (n_2820));
  NA2X1 g62403(.A (n_2427), .B (n_2428), .Q (n_2819));
  NA2X1 g62404(.A (n_2403), .B (n_2406), .Q (n_2818));
  AN211X1 g62405(.A (n_2164), .B (n_4965), .C (n_2341), .D (n_2340), .Q
       (n_2817));
  NA2X1 g62406(.A (n_2450), .B (n_2447), .Q (n_2816));
  NA2X1 g62407(.A (n_2445), .B (n_2446), .Q (n_2815));
  AN211X1 g62408(.A (n_2164), .B (n_4934), .C (n_2337), .D (n_2338), .Q
       (n_2814));
  NA2X1 g62409(.A (n_2474), .B (n_2336), .Q (n_2813));
  AN221X1 g62410(.A (n_4951), .B (n_2173), .C (n_4950), .D (n_1600), .E
       (n_2423), .Q (n_2812));
  AN221X1 g62411(.A (n_4978), .B (n_2171), .C (n_4977), .D (n_2167), .E
       (n_2422), .Q (n_2811));
  AN211X1 g62416(.A (n_2164), .B (n_4903), .C (n_2329), .D (n_2330), .Q
       (n_2807));
  NA2X1 g62417(.A (n_2451), .B (n_2311), .Q (n_2806));
  NA2X2 g62418(.A (n_2400), .B (n_2409), .Q (n_2805));
  NA2X1 g62419(.A (n_2413), .B (n_2391), .Q (n_2804));
  NA2X1 g62420(.A (n_2404), .B (n_2387), .Q (n_2803));
  NA2X1 g62422(.A (n_2419), .B (n_2418), .Q (n_2802));
  NA2X1 g62426(.A (n_2420), .B (n_6753), .Q (n_2800));
  NA2X1 g62428(.A (n_2407), .B (n_2408), .Q (n_2798));
  NA3X1 g62429(.A (n_2250), .B (n_2370), .C (n_2075), .Q
       (csr_data_out[9]));
  NA3X1 g62430(.A (n_2248), .B (n_2331), .C (n_2033), .Q
       (csr_data_out[5]));
  NA6X1 g62431(.A (n_2036), .B (n_2030), .C (n_2125), .D (n_2123), .E
       (n_2001), .F (n_2025), .Q (csr_data_out[2]));
  NA6X1 g62432(.A (n_2133), .B (n_2275), .C (n_2028), .D (n_2031), .E
       (n_2121), .F (n_2119), .Q (csr_data_out[3]));
  NA3X1 g62433(.A (n_2249), .B (n_2359), .C (n_2041), .Q
       (csr_data_out[6]));
  NA6X1 g62434(.A (n_2053), .B (n_2044), .C (n_2132), .D (n_2134), .E
       (n_2006), .F (n_2029), .Q (csr_data_out[8]));
  NA6X1 g62435(.A (n_2038), .B (n_2032), .C (n_2126), .D (n_2127), .E
       (n_2002), .F (n_2026), .Q (csr_data_out[4]));
  OR2X1 g62436(.A (n_2321), .B (n_2589), .Q (n_2886));
  NO2X1 g62437(.A (n_2321), .B (n_2586), .Q (n_2884));
  OR2X1 g62438(.A (n_2321), .B (n_2588), .Q (n_2883));
  NO2X1 g62439(.A (n_2321), .B (n_2587), .Q (n_2881));
  INX1 g62440(.A (n_2796), .Q (n_2797));
  AN22X1 g62441(.A (n_2185), .B (n_4552), .C (n_2187), .D (n_4551), .Q
       (n_2793));
  NA3X1 g62442(.A (n_2381), .B (n_2262), .C (n_1906), .Q (n_2792));
  AN22X1 g62443(.A (n_2171), .B (n_4575), .C (n_2167), .D (n_4574), .Q
       (n_2791));
  AN22X1 g62444(.A (n_1596), .B (n_5421), .C (n_2188), .D (n_5418), .Q
       (n_2790));
  AN22X1 g62445(.A (n_1595), .B (n_5452), .C (n_2188), .D (n_5449), .Q
       (n_2789));
  AN22X1 g62446(.A (n_1595), .B (n_4677), .C (n_2188), .D (n_4674), .Q
       (n_2788));
  AO22X1 g62448(.A (n_1595), .B (n_5173), .C (n_2188), .D (n_5170), .Q
       (n_2786));
  AN22X1 g62449(.A (n_2185), .B (n_4583), .C (n_2187), .D (n_4582), .Q
       (n_2785));
  AN22X1 g62450(.A (n_2185), .B (n_4831), .C (n_2187), .D (n_4830), .Q
       (n_2784));
  AN22X1 g62451(.A (n_2185), .B (n_5110), .C (n_2187), .D (n_5109), .Q
       (n_2783));
  AN22X1 g62452(.A (n_2185), .B (n_4707), .C (n_2187), .D (n_4706), .Q
       (n_2782));
  AN22X1 g62453(.A (n_2185), .B (n_4676), .C (n_2187), .D (n_4675), .Q
       (n_2781));
  AN22X1 g62454(.A (n_2185), .B (n_4645), .C (n_2187), .D (n_4644), .Q
       (n_2780));
  AN22X1 g62455(.A (n_2185), .B (n_5172), .C (n_2187), .D (n_5171), .Q
       (n_2779));
  AN22X1 g62456(.A (n_2185), .B (n_4614), .C (n_2187), .D (n_4613), .Q
       (n_2778));
  AN22X1 g62457(.A (n_1596), .B (n_4832), .C (n_2188), .D (n_4829), .Q
       (n_2777));
  AN22X1 g62458(.A (n_2202), .B (n_4834), .C (n_2198), .D (n_4833), .Q
       (n_2776));
  AN22X1 g62459(.A (n_2202), .B (n_5113), .C (n_2198), .D (n_5112), .Q
       (n_2775));
  AN22X1 g62460(.A (n_1595), .B (n_5514), .C (n_2188), .D (n_5511), .Q
       (n_2774));
  AO22X1 g62461(.A (n_2202), .B (n_5454), .C (n_2198), .D (n_5453), .Q
       (n_2773));
  AN22X1 g62462(.A (n_2202), .B (n_4710), .C (n_2198), .D (n_4709), .Q
       (n_2772));
  AO22X1 g62463(.A (n_2202), .B (n_5516), .C (n_2198), .D (n_5515), .Q
       (n_2771));
  AN22X1 g62464(.A (n_2202), .B (n_4679), .C (n_2198), .D (n_4678), .Q
       (n_2770));
  AO22X1 g62465(.A (n_2202), .B (n_5361), .C (n_2198), .D (n_5360), .Q
       (n_2769));
  AN22X1 g62466(.A (n_2202), .B (n_4648), .C (n_2198), .D (n_4647), .Q
       (n_2768));
  AN22X1 g62467(.A (n_2202), .B (n_5175), .C (n_2198), .D (n_5174), .Q
       (n_2767));
  AO22X1 g62469(.A (n_2202), .B (n_5423), .C (n_2198), .D (n_5422), .Q
       (n_2765));
  AN22X1 g62470(.A (n_2200), .B (n_4587), .C (n_2153), .D (n_4589), .Q
       (n_2764));
  AN22X1 g62471(.A (n_2200), .B (n_4835), .C (n_2153), .D (n_4837), .Q
       (n_2763));
  AN22X1 g62472(.A (n_2200), .B (n_4680), .C (n_2153), .D (n_4682), .Q
       (n_2762));
  AN22X1 g62473(.A (n_2200), .B (n_4649), .C (n_2153), .D (n_4651), .Q
       (n_2761));
  AN22X1 g62474(.A (n_2200), .B (n_5176), .C (n_2153), .D (n_5178), .Q
       (n_2760));
  AN22X1 g62475(.A (n_2200), .B (n_4618), .C (n_2153), .D (n_4620), .Q
       (n_2759));
  AN22X1 g62476(.A (n_2193), .B (n_5437), .C (n_2195), .D (n_5438), .Q
       (n_2758));
  AO22X1 g62477(.A (n_2196), .B (n_5439), .C (n_2181), .D (n_5433), .Q
       (n_2757));
  AN22X1 g62478(.A (n_2191), .B (n_5440), .C (n_2183), .D (n_5436), .Q
       (n_2756));
  AN22X1 g62479(.A (n_2154), .B (n_5432), .C (n_2156), .D (n_5431), .Q
       (n_2755));
  AO22X1 g62480(.A (n_2150), .B (n_5428), .C (n_2152), .D (n_5427), .Q
       (n_2754));
  AN22X1 g62481(.A (n_2196), .B (n_5129), .C (n_2195), .D (n_5128), .Q
       (n_2753));
  AO22X1 g62482(.A (n_2196), .B (n_5470), .C (n_2195), .D (n_5469), .Q
       (n_2752));
  AN22X1 g62483(.A (n_2193), .B (n_4693), .C (n_2195), .D (n_4694), .Q
       (n_2751));
  AO22X1 g62484(.A (n_2193), .B (n_5530), .C (n_2195), .D (n_5531), .Q
       (n_2750));
  AN22X1 g62485(.A (n_2193), .B (n_4662), .C (n_2195), .D (n_4663), .Q
       (n_2749));
  AO22X1 g62486(.A (n_2196), .B (n_5191), .C (n_2195), .D (n_5190), .Q
       (n_2748));
  AN22X1 g62487(.A (n_2181), .B (n_5123), .C (n_2179), .D (n_5125), .Q
       (n_2747));
  AN22X1 g62488(.A (n_2181), .B (n_5464), .C (n_2177), .D (n_5465), .Q
       (n_2746));
  AN22X1 g62489(.A (n_2179), .B (n_4691), .C (n_2177), .D (n_4690), .Q
       (n_2745));
  AN22X1 g62490(.A (n_2181), .B (n_4658), .C (n_2179), .D (n_4660), .Q
       (n_2744));
  AN22X1 g62491(.A (n_2191), .B (n_5130), .C (n_2183), .D (n_5126), .Q
       (n_2743));
  AN22X1 g62492(.A (n_2193), .B (n_5127), .C (n_2177), .D (n_5124), .Q
       (n_2742));
  AN22X1 g62493(.A (n_2193), .B (n_5468), .C (n_2179), .D (n_5466), .Q
       (n_2741));
  AO22X1 g62494(.A (n_2196), .B (n_5532), .C (n_2177), .D (n_5527), .Q
       (n_2740));
  AN22X1 g62495(.A (n_2196), .B (n_4695), .C (n_2181), .D (n_4689), .Q
       (n_2739));
  AN22X1 g62496(.A (n_2191), .B (n_4696), .C (n_2183), .D (n_4692), .Q
       (n_2738));
  AN22X1 g62497(.A (n_2196), .B (n_4664), .C (n_2177), .D (n_4659), .Q
       (n_2737));
  AN22X1 g62498(.A (n_2191), .B (n_4665), .C (n_2183), .D (n_4661), .Q
       (n_2736));
  AO22X1 g62499(.A (n_2193), .B (n_5189), .C (n_2179), .D (n_5187), .Q
       (n_2735));
  AO22X1 g62500(.A (n_2150), .B (n_4591), .C (n_2152), .D (n_4590), .Q
       (n_2734));
  AN22X1 g62501(.A (n_2154), .B (n_4843), .C (n_2156), .D (n_4842), .Q
       (n_2733));
  AN22X1 g62502(.A (n_2150), .B (n_4839), .C (n_2152), .D (n_4838), .Q
       (n_2732));
  AO22X1 g62503(.A (n_2154), .B (n_5122), .C (n_2156), .D (n_5121), .Q
       (n_2731));
  AO22X1 g62504(.A (n_2150), .B (n_5118), .C (n_2152), .D (n_5117), .Q
       (n_2730));
  AN22X1 g62505(.A (n_2154), .B (n_5525), .C (n_2156), .D (n_5524), .Q
       (n_2729));
  AN22X1 g62506(.A (n_2154), .B (n_5463), .C (n_2156), .D (n_5462), .Q
       (n_2728));
  AO22X1 g62507(.A (n_2150), .B (n_5459), .C (n_2152), .D (n_5458), .Q
       (n_2727));
  AN22X1 g62508(.A (n_2154), .B (n_4719), .C (n_2160), .D (n_4712), .Q
       (n_2726));
  AO22X1 g62509(.A (n_2150), .B (n_4715), .C (n_2152), .D (n_4714), .Q
       (n_2725));
  AN22X1 g62511(.A (n_2154), .B (n_4688), .C (n_2156), .D (n_4687), .Q
       (n_2723));
  AN22X1 g62512(.A (n_2150), .B (n_4684), .C (n_2152), .D (n_4683), .Q
       (n_2722));
  AO22X1 g62513(.A (n_2154), .B (n_5370), .C (n_2156), .D (n_5369), .Q
       (n_2721));
  AO22X1 g62514(.A (n_2150), .B (n_5366), .C (n_2152), .D (n_5365), .Q
       (n_2720));
  AO22X1 g62515(.A (n_2154), .B (n_4657), .C (n_2156), .D (n_4656), .Q
       (n_2719));
  AN22X1 g62517(.A (n_2150), .B (n_4653), .C (n_2152), .D (n_4652), .Q
       (n_2717));
  AO22X1 g62518(.A (n_2154), .B (n_4626), .C (n_2156), .D (n_4625), .Q
       (n_2716));
  AN22X1 g62519(.A (n_2150), .B (n_5180), .C (n_2152), .D (n_5179), .Q
       (n_2715));
  AO22X1 g62520(.A (n_2150), .B (n_4622), .C (n_2152), .D (n_4621), .Q
       (n_2714));
  AO22X1 g62521(.A (n_2150), .B (n_5521), .C (n_2152), .D (n_5520), .Q
       (n_2713));
  AN22X1 g62522(.A (n_2173), .B (n_5447), .C (n_2169), .D (n_5441), .Q
       (n_2712));
  AN22X1 g62523(.A (n_2165), .B (n_5445), .C (n_1600), .D (n_5446), .Q
       (n_2711));
  AN22X1 g62524(.A (n_2185), .B (n_5079), .C (n_2187), .D (n_5078), .Q
       (n_2710));
  AN22X1 g62525(.A (n_2185), .B (n_5048), .C (n_2187), .D (n_5047), .Q
       (n_2709));
  AN22X1 g62526(.A (n_2185), .B (n_5234), .C (n_2187), .D (n_5233), .Q
       (n_2708));
  AN22X1 g62527(.A (n_1596), .B (n_5080), .C (n_2188), .D (n_5077), .Q
       (n_2707));
  AN22X1 g62528(.A (n_2202), .B (n_5082), .C (n_2198), .D (n_5081), .Q
       (n_2706));
  AN22X1 g62529(.A (n_2200), .B (n_5083), .C (n_2153), .D (n_5085), .Q
       (n_2705));
  AN22X1 g62530(.A (n_2202), .B (n_5051), .C (n_2198), .D (n_5050), .Q
       (n_2704));
  AN22X1 g62531(.A (n_2200), .B (n_5052), .C (n_2153), .D (n_5054), .Q
       (n_2703));
  AN22X1 g62532(.A (n_1596), .B (n_5390), .C (n_2188), .D (n_5387), .Q
       (n_2702));
  AO22X1 g62533(.A (n_2202), .B (n_5392), .C (n_2198), .D (n_5391), .Q
       (n_2701));
  AN22X1 g62534(.A (n_1595), .B (n_5266), .C (n_2188), .D (n_5263), .Q
       (n_2700));
  AO22X1 g62535(.A (n_2202), .B (n_5268), .C (n_2198), .D (n_5267), .Q
       (n_2699));
  AN22X1 g62536(.A (n_2200), .B (n_5269), .C (n_2153), .D (n_5271), .Q
       (n_2698));
  AN22X1 g62537(.A (n_1596), .B (n_5235), .C (n_2188), .D (n_5232), .Q
       (n_2697));
  AN22X1 g62538(.A (n_2202), .B (n_5237), .C (n_2198), .D (n_5236), .Q
       (n_2696));
  AN22X1 g62539(.A (n_2200), .B (n_5238), .C (n_2153), .D (n_5240), .Q
       (n_2695));
  AN22X1 g62540(.A (n_2200), .B (n_5486), .C (n_2153), .D (n_5488), .Q
       (n_2694));
  AN22X1 g62541(.A (n_2200), .B (n_4556), .C (n_2153), .D (n_4558), .Q
       (n_2693));
  AN22X1 g62542(.A (n_2185), .B (n_5482), .C (n_2187), .D (n_5481), .Q
       (n_2692));
  OR2X1 g62543(.A (n_2380), .B (n_2382), .Q (n_2691));
  AN22X1 g62544(.A (n_2179), .B (n_4598), .C (n_2177), .D (n_4597), .Q
       (n_2690));
  AN22X1 g62545(.A (n_2179), .B (n_4846), .C (n_2177), .D (n_4845), .Q
       (n_2689));
  AN22X1 g62546(.A (n_2179), .B (n_5094), .C (n_2177), .D (n_5093), .Q
       (n_2688));
  AN22X1 g62547(.A (n_2181), .B (n_5061), .C (n_2177), .D (n_5062), .Q
       (n_2687));
  AN22X1 g62548(.A (n_2179), .B (n_4722), .C (n_2177), .D (n_4721), .Q
       (n_2686));
  AN22X1 g62549(.A (n_2179), .B (n_5373), .C (n_2177), .D (n_5372), .Q
       (n_2685));
  AN22X1 g62550(.A (n_2181), .B (n_5371), .C (n_2195), .D (n_5376), .Q
       (n_2684));
  AN22X1 g62551(.A (n_2179), .B (n_4629), .C (n_2177), .D (n_4628), .Q
       (n_2683));
  AN22X1 g62552(.A (n_2169), .B (n_5131), .C (n_2171), .D (n_5133), .Q
       (n_2682));
  AN22X1 g62553(.A (n_2165), .B (n_5135), .C (n_1600), .D (n_5136), .Q
       (n_2681));
  AN22X1 g62554(.A (n_2173), .B (n_5478), .C (n_2169), .D (n_5472), .Q
       (n_2680));
  AN22X1 g62555(.A (n_2165), .B (n_5476), .C (n_1600), .D (n_5477), .Q
       (n_2679));
  AN22X1 g62556(.A (n_2169), .B (n_5534), .C (n_2171), .D (n_5536), .Q
       (n_2678));
  AN22X1 g62557(.A (n_2202), .B (n_5485), .C (n_2198), .D (n_5484), .Q
       (n_2677));
  AN22X1 g62558(.A (n_2165), .B (n_5538), .C (n_2167), .D (n_5535), .Q
       (n_2676));
  AN22X1 g62559(.A (n_1595), .B (n_4553), .C (n_2188), .D (n_4550), .Q
       (n_2675));
  AN22X1 g62560(.A (n_1595), .B (n_5483), .C (n_2188), .D (n_5480), .Q
       (n_2674));
  AN22X1 g62561(.A (n_2202), .B (n_4555), .C (n_2198), .D (n_4554), .Q
       (n_2673));
  AN22X1 g62562(.A (n_2165), .B (n_4701), .C (n_1600), .D (n_4702), .Q
       (n_2672));
  AN22X1 g62563(.A (n_2171), .B (n_4699), .C (n_2167), .D (n_4698), .Q
       (n_2671));
  AN22X1 g62564(.A (n_2173), .B (n_4703), .C (n_2169), .D (n_4697), .Q
       (n_2670));
  AN22X1 g62565(.A (n_2171), .B (n_4668), .C (n_2167), .D (n_4667), .Q
       (n_2669));
  AN22X1 g62566(.A (n_2173), .B (n_4672), .C (n_2169), .D (n_4666), .Q
       (n_2668));
  AN22X1 g62567(.A (n_2165), .B (n_4670), .C (n_1600), .D (n_4671), .Q
       (n_2667));
  AO22X1 g62568(.A (n_2169), .B (n_5193), .C (n_2171), .D (n_5195), .Q
       (n_2666));
  AN22X1 g62569(.A (n_2191), .B (n_4603), .C (n_2183), .D (n_4599), .Q
       (n_2665));
  AN22X1 g62570(.A (n_2196), .B (n_4602), .C (n_2181), .D (n_4596), .Q
       (n_2664));
  AN22X1 g62571(.A (n_2193), .B (n_4600), .C (n_2195), .D (n_4601), .Q
       (n_2663));
  AN22X1 g62572(.A (n_2191), .B (n_4851), .C (n_2183), .D (n_4847), .Q
       (n_2662));
  AN22X1 g62573(.A (n_2196), .B (n_4850), .C (n_2181), .D (n_4844), .Q
       (n_2661));
  AN22X1 g62574(.A (n_2193), .B (n_4848), .C (n_2195), .D (n_4849), .Q
       (n_2660));
  AN22X1 g62575(.A (n_2191), .B (n_5099), .C (n_2183), .D (n_5095), .Q
       (n_2659));
  AN22X1 g62576(.A (n_2196), .B (n_5098), .C (n_2181), .D (n_5092), .Q
       (n_2658));
  AN22X1 g62577(.A (n_2193), .B (n_5096), .C (n_2195), .D (n_5097), .Q
       (n_2657));
  AN22X1 g62578(.A (n_2196), .B (n_5067), .C (n_2195), .D (n_5066), .Q
       (n_2656));
  AN22X1 g62579(.A (n_2191), .B (n_5068), .C (n_2183), .D (n_5064), .Q
       (n_2655));
  AN22X1 g62580(.A (n_2193), .B (n_5065), .C (n_2179), .D (n_5063), .Q
       (n_2654));
  AN22X1 g62581(.A (n_2191), .B (n_4727), .C (n_2183), .D (n_4723), .Q
       (n_2653));
  AO22X1 g62582(.A (n_2193), .B (n_4724), .C (n_2196), .D (n_4726), .Q
       (n_2652));
  AO22X1 g62583(.A (n_2191), .B (n_5409), .C (n_2183), .D (n_5405), .Q
       (n_2651));
  AO22X1 g62584(.A (n_2196), .B (n_5408), .C (n_2181), .D (n_5402), .Q
       (n_2650));
  AN22X1 g62585(.A (n_2191), .B (n_5378), .C (n_2183), .D (n_5374), .Q
       (n_2649));
  AN22X1 g62586(.A (n_2193), .B (n_5375), .C (n_2196), .D (n_5377), .Q
       (n_2648));
  AN22X1 g62587(.A (n_2191), .B (n_4634), .C (n_2183), .D (n_4630), .Q
       (n_2647));
  AN22X1 g62588(.A (n_2196), .B (n_4633), .C (n_2181), .D (n_4627), .Q
       (n_2646));
  AN22X1 g62589(.A (n_2193), .B (n_4631), .C (n_2195), .D (n_4632), .Q
       (n_2645));
  AN22X1 g62590(.A (n_2179), .B (n_5249), .C (n_2177), .D (n_5248), .Q
       (n_2644));
  AN22X1 g62591(.A (n_2181), .B (n_5247), .C (n_2195), .D (n_5252), .Q
       (n_2643));
  AN22X1 g62592(.A (n_2181), .B (n_5495), .C (n_2177), .D (n_5496), .Q
       (n_2642));
  AN22X1 g62593(.A (n_2179), .B (n_4567), .C (n_2177), .D (n_4566), .Q
       (n_2641));
  AN22X1 g62594(.A (n_2179), .B (n_5280), .C (n_2177), .D (n_5279), .Q
       (n_2640));
  AN22X1 g62595(.A (n_2181), .B (n_5278), .C (n_2195), .D (n_5283), .Q
       (n_2639));
  AN22X1 g62596(.A (n_2191), .B (n_5254), .C (n_2183), .D (n_5250), .Q
       (n_2638));
  AN22X1 g62597(.A (n_2193), .B (n_5251), .C (n_2196), .D (n_5253), .Q
       (n_2637));
  AN22X1 g62598(.A (n_2154), .B (n_5494), .C (n_2156), .D (n_5493), .Q
       (n_2636));
  AN22X1 g62599(.A (n_2150), .B (n_5490), .C (n_2152), .D (n_5489), .Q
       (n_2635));
  AN22X1 g62600(.A (n_2196), .B (n_5501), .C (n_2195), .D (n_5500), .Q
       (n_2634));
  AN22X1 g62601(.A (n_2191), .B (n_5502), .C (n_2183), .D (n_5498), .Q
       (n_2633));
  AN22X1 g62602(.A (n_2193), .B (n_5499), .C (n_2179), .D (n_5497), .Q
       (n_2632));
  AN22X1 g62603(.A (n_2150), .B (n_4560), .C (n_2152), .D (n_4559), .Q
       (n_2631));
  AN22X1 g62604(.A (n_2191), .B (n_4572), .C (n_2183), .D (n_4568), .Q
       (n_2630));
  AN22X1 g62605(.A (n_2196), .B (n_4571), .C (n_2181), .D (n_4565), .Q
       (n_2629));
  AN22X1 g62606(.A (n_2193), .B (n_4569), .C (n_2195), .D (n_4570), .Q
       (n_2628));
  AN22X1 g62607(.A (n_2191), .B (n_5285), .C (n_2183), .D (n_5281), .Q
       (n_2627));
  AN22X1 g62608(.A (n_2193), .B (n_5282), .C (n_2196), .D (n_5284), .Q
       (n_2626));
  AN22X1 g62609(.A (n_2154), .B (n_4564), .C (n_2156), .D (n_4563), .Q
       (n_2625));
  AN22X1 g62610(.A (n_2154), .B (n_5091), .C (n_2156), .D (n_5090), .Q
       (n_2624));
  AN22X1 g62611(.A (n_2150), .B (n_5087), .C (n_2152), .D (n_5086), .Q
       (n_2623));
  AN22X1 g62612(.A (n_2154), .B (n_5060), .C (n_2160), .D (n_5053), .Q
       (n_2622));
  AN22X1 g62613(.A (n_2150), .B (n_5056), .C (n_2152), .D (n_5055), .Q
       (n_2621));
  AN22X1 g62614(.A (n_2154), .B (n_5401), .C (n_2156), .D (n_5400), .Q
       (n_2620));
  AO22X1 g62615(.A (n_2150), .B (n_5397), .C (n_2152), .D (n_5396), .Q
       (n_2619));
  AN22X1 g62617(.A (n_2154), .B (n_5277), .C (n_2156), .D (n_5276), .Q
       (n_2617));
  AN22X1 g62618(.A (n_2150), .B (n_5273), .C (n_2152), .D (n_5272), .Q
       (n_2616));
  AN22X1 g62619(.A (n_2154), .B (n_5246), .C (n_2156), .D (n_5245), .Q
       (n_2615));
  AN22X1 g62620(.A (n_2150), .B (n_5242), .C (n_2152), .D (n_5241), .Q
       (n_2614));
  AN22X1 g62621(.A (n_2156), .B (n_5059), .C (n_2164), .D (n_5058), .Q
       (n_2613));
  AN22X1 g62622(.A (n_2156), .B (n_4718), .C (n_2164), .D (n_4717), .Q
       (n_2612));
  AO22X1 g62623(.A (n_2156), .B (n_4594), .C (n_2164), .D (n_4593), .Q
       (n_2611));
  AN22X1 g62624(.A (n_2173), .B (n_4610), .C (n_1598), .D (n_4609), .Q
       (n_2610));
  AN22X1 g62625(.A (n_2169), .B (n_5410), .C (n_2171), .D (n_5412), .Q
       (n_2609));
  AN22X1 g62626(.A (n_2165), .B (n_4608), .C (n_2171), .D (n_4606), .Q
       (n_2608));
  AO22X1 g62627(.A (n_2173), .B (n_4858), .C (n_2169), .D (n_4852), .Q
       (n_2607));
  AN22X1 g62628(.A (n_2169), .B (n_5100), .C (n_2171), .D (n_5102), .Q
       (n_2606));
  AN22X1 g62629(.A (n_2165), .B (n_5104), .C (n_2167), .D (n_5101), .Q
       (n_2605));
  AN22X1 g62631(.A (n_2169), .B (n_5069), .C (n_2167), .D (n_5070), .Q
       (n_2603));
  AN22X1 g62632(.A (n_2165), .B (n_5073), .C (n_2171), .D (n_5071), .Q
       (n_2602));
  AN22X1 g62633(.A (n_2169), .B (n_4728), .C (n_2167), .D (n_4729), .Q
       (n_2601));
  AN22X1 g62634(.A (n_1598), .B (n_4733), .C (n_2171), .D (n_4730), .Q
       (n_2600));
  AN22X1 g62635(.A (n_2165), .B (n_4732), .C (n_2173), .D (n_4734), .Q
       (n_2599));
  AN22X1 g62636(.A (n_2173), .B (n_5385), .C (n_2169), .D (n_5379), .Q
       (n_2598));
  AN22X1 g62637(.A (n_2165), .B (n_5383), .C (n_1600), .D (n_5384), .Q
       (n_2597));
  AN22X1 g62638(.A (n_2165), .B (n_5414), .C (n_2167), .D (n_5411), .Q
       (n_2596));
  AN22X1 g62639(.A (n_2173), .B (n_4641), .C (n_2171), .D (n_4637), .Q
       (n_2595));
  AN22X1 g62640(.A (n_2165), .B (n_4639), .C (n_1598), .D (n_4640), .Q
       (n_2594));
  AN22X1 g62641(.A (n_2173), .B (n_5509), .C (n_2171), .D (n_5505), .Q
       (n_2593));
  AN22X1 g62642(.A (n_2169), .B (n_5503), .C (n_2167), .D (n_5504), .Q
       (n_2592));
  AN22X1 g62643(.A (n_2165), .B (n_5507), .C (n_1598), .D (n_5508), .Q
       (n_2591));
  AN22X1 g62644(.A (n_2264), .B (n_1727), .C (n_5604), .D (n_5606), .Q
       (n_2796));
  AO21X1 g62645(.A (n_6461), .B (n_1840), .C (n_2380), .Q (n_2795));
  ON21X1 g62646(.A (n_6065), .B (n_1841), .C (n_2262), .Q (n_2794));
  AN22X1 g62647(.A (n_2200), .B (n_4928), .C (n_2153), .D (n_4930), .Q
       (n_2585));
  AN22X1 g62648(.A (n_2165), .B (n_4577), .C (n_1598), .D (n_4578), .Q
       (n_2584));
  AN22X1 g62649(.A (n_2173), .B (n_5292), .C (n_1598), .D (n_5291), .Q
       (n_2583));
  AN22X1 g62650(.A (n_2169), .B (n_5286), .C (n_2167), .D (n_5287), .Q
       (n_2582));
  AN22X1 g62651(.A (n_2165), .B (n_5290), .C (n_2171), .D (n_5288), .Q
       (n_2581));
  AN22X1 g62652(.A (n_2169), .B (n_5255), .C (n_2167), .D (n_5256), .Q
       (n_2580));
  AN22X1 g62653(.A (n_2173), .B (n_5261), .C (n_2171), .D (n_5257), .Q
       (n_2579));
  AN22X1 g62654(.A (n_2202), .B (n_5206), .C (n_2198), .D (n_5205), .Q
       (n_2578));
  AN22X1 g62655(.A (n_2202), .B (n_5144), .C (n_2198), .D (n_5143), .Q
       (n_2577));
  AN22X1 g62656(.A (n_2202), .B (n_5020), .C (n_2198), .D (n_5019), .Q
       (n_2576));
  AO22X1 g62657(.A (n_2202), .B (n_5330), .C (n_2198), .D (n_5329), .Q
       (n_2575));
  AO22X1 g62658(.A (n_2202), .B (n_5299), .C (n_2198), .D (n_5298), .Q
       (n_2574));
  AN22X1 g62660(.A (n_2185), .B (n_5203), .C (n_2187), .D (n_5202), .Q
       (n_2572));
  NO2X1 g62661(.A (n_2354), .B (n_2356), .Q (n_2571));
  AN22X1 g62662(.A (n_2185), .B (n_5141), .C (n_2187), .D (n_5140), .Q
       (n_2570));
  NO2X1 g62663(.A (n_2353), .B (n_2355), .Q (n_2569));
  AN22X1 g62664(.A (n_2185), .B (n_5017), .C (n_2187), .D (n_5016), .Q
       (n_2568));
  AN22X1 g62665(.A (n_1596), .B (n_5297), .C (n_2188), .D (n_5294), .Q
       (n_2567));
  AN22X1 g62668(.A (n_2181), .B (n_5030), .C (n_2177), .D (n_5031), .Q
       (n_2564));
  AN22X1 g62669(.A (n_2181), .B (n_5340), .C (n_2177), .D (n_5341), .Q
       (n_2563));
  AO22X1 g62671(.A (n_2191), .B (n_5223), .C (n_2183), .D (n_5219), .Q
       (n_2561));
  AO22X1 g62672(.A (n_2193), .B (n_5220), .C (n_2195), .D (n_5221), .Q
       (n_2560));
  AO22X1 g62674(.A (n_2191), .B (n_5161), .C (n_2183), .D (n_5157), .Q
       (n_2558));
  AO22X1 g62675(.A (n_2193), .B (n_5158), .C (n_2179), .D (n_5156), .Q
       (n_2557));
  AN22X1 g62676(.A (n_2196), .B (n_5036), .C (n_2195), .D (n_5035), .Q
       (n_2556));
  AN22X1 g62677(.A (n_2191), .B (n_5037), .C (n_2183), .D (n_5033), .Q
       (n_2555));
  AN22X1 g62678(.A (n_2193), .B (n_5034), .C (n_2179), .D (n_5032), .Q
       (n_2554));
  AN22X1 g62679(.A (n_2196), .B (n_5346), .C (n_2179), .D (n_5342), .Q
       (n_2553));
  AN22X1 g62680(.A (n_2191), .B (n_5347), .C (n_2183), .D (n_5343), .Q
       (n_2552));
  AN22X1 g62681(.A (n_2193), .B (n_5344), .C (n_2195), .D (n_5345), .Q
       (n_2551));
  AO22X1 g62682(.A (n_2191), .B (n_5316), .C (n_2183), .D (n_5312), .Q
       (n_2550));
  AO22X1 g62683(.A (n_2193), .B (n_5313), .C (n_2179), .D (n_5311), .Q
       (n_2549));
  AN22X1 g62684(.A (n_2200), .B (n_5207), .C (n_2153), .D (n_5209), .Q
       (n_2548));
  AN22X1 g62685(.A (n_2200), .B (n_5145), .C (n_2153), .D (n_5147), .Q
       (n_2547));
  AN22X1 g62687(.A (n_2200), .B (n_5331), .C (n_2153), .D (n_5333), .Q
       (n_2545));
  AN22X1 g62688(.A (n_2200), .B (n_5300), .C (n_2153), .D (n_5302), .Q
       (n_2544));
  AO22X1 g62689(.A (n_2176), .B (n_5444), .C (n_1813), .D (n_5448), .Q
       (n_2543));
  NO2X1 g62691(.A (n_2347), .B (n_2348), .Q (n_2541));
  AN22X1 g62692(.A (n_2150), .B (n_5211), .C (n_2152), .D (n_5210), .Q
       (n_2540));
  AN22X1 g62695(.A (n_2150), .B (n_5149), .C (n_2152), .D (n_5148), .Q
       (n_2537));
  NO2X1 g62696(.A (n_2345), .B (n_2346), .Q (n_2536));
  AN22X1 g62697(.A (n_2154), .B (n_5029), .C (n_2156), .D (n_5028), .Q
       (n_2535));
  AO22X1 g62698(.A (n_2150), .B (n_5025), .C (n_2152), .D (n_5024), .Q
       (n_2534));
  AO22X1 g62699(.A (n_2154), .B (n_5339), .C (n_2156), .D (n_5338), .Q
       (n_2533));
  AN22X1 g62700(.A (n_2150), .B (n_5335), .C (n_2152), .D (n_5334), .Q
       (n_2532));
  AN22X1 g62701(.A (n_2154), .B (n_5308), .C (n_2156), .D (n_5307), .Q
       (n_2531));
  AN22X1 g62702(.A (n_2150), .B (n_5304), .C (n_2152), .D (n_5303), .Q
       (n_2530));
  AN22X1 g62703(.A (n_2202), .B (n_4958), .C (n_2198), .D (n_4957), .Q
       (n_2529));
  AN22X1 g62704(.A (n_1595), .B (n_4956), .C (n_2188), .D (n_4953), .Q
       (n_2528));
  AN22X1 g62705(.A (n_2185), .B (n_4955), .C (n_2187), .D (n_4954), .Q
       (n_2527));
  ON22X1 g62706(.A (n_2201), .B (n_1677), .C (n_1573), .D (n_1676), .Q
       (n_2526));
  ON21X1 g62707(.A (n_1601), .B (n_1678), .C (n_1870), .Q (n_2525));
  ON21X1 g62708(.A (n_1601), .B (n_1668), .C (n_1868), .Q (n_2524));
  ON21X1 g62709(.A (n_1601), .B (n_1675), .C (n_1867), .Q (n_2523));
  AN21X1 g62710(.A (n_2176), .B (n_4700), .C (n_1869), .Q (n_2522));
  AN22X1 g62711(.A (n_2176), .B (n_4669), .C (n_1813), .D (n_4673), .Q
       (n_2521));
  AO22X1 g62712(.A (n_2176), .B (n_5196), .C (n_1813), .D (n_5200), .Q
       (n_2520));
  AN22X1 g62713(.A (n_2154), .B (n_4967), .C (n_2156), .D (n_4966), .Q
       (n_2519));
  AN22X1 g62715(.A (n_2185), .B (n_4986), .C (n_2187), .D (n_4985), .Q
       (n_2517));
  AN22X1 g62716(.A (n_1595), .B (n_4925), .C (n_2188), .D (n_4922), .Q
       (n_2516));
  AO22X1 g62717(.A (n_2202), .B (n_4927), .C (n_2198), .D (n_4926), .Q
       (n_2515));
  AN21X1 g62718(.A (n_2188), .B (n_4984), .C (n_2332), .Q (n_2514));
  AN22X1 g62719(.A (n_2202), .B (n_4989), .C (n_2198), .D (n_4988), .Q
       (n_2513));
  ON21X1 g62720(.A (n_1601), .B (n_1674), .C (n_1866), .Q (n_2512));
  NO2X1 g62721(.A (n_2326), .B (n_2327), .Q (n_2511));
  NO2X1 g62722(.A (n_2324), .B (n_2325), .Q (n_2510));
  NO2X1 g62723(.A (n_2377), .B (n_2376), .Q (n_2509));
  AN22X1 g62724(.A (n_2169), .B (n_5162), .C (n_2167), .D (n_5163), .Q
       (n_2508));
  NO2X1 g62725(.A (n_2320), .B (n_2378), .Q (n_2507));
  AN22X1 g62726(.A (n_2165), .B (n_5166), .C (n_1600), .D (n_5167), .Q
       (n_2506));
  AO22X1 g62727(.A (n_2176), .B (n_4855), .C (n_1813), .D (n_4859), .Q
       (n_2505));
  ON21X1 g62728(.A (n_1601), .B (n_1670), .C (n_1865), .Q (n_2504));
  ON22X1 g62729(.A (n_1601), .B (n_1683), .C (n_1812), .D (n_1710), .Q
       (n_2503));
  AN22X1 g62730(.A (n_2173), .B (n_5044), .C (n_1600), .D (n_5043), .Q
       (n_2502));
  AN22X1 g62731(.A (n_2169), .B (n_5038), .C (n_2167), .D (n_5039), .Q
       (n_2501));
  AN22X1 g62732(.A (n_2165), .B (n_5042), .C (n_2171), .D (n_5040), .Q
       (n_2500));
  AN22X1 g62733(.A (n_2176), .B (n_4731), .C (n_1813), .D (n_4735), .Q
       (n_2499));
  ON21X1 g62734(.A (n_1601), .B (n_1666), .C (n_1863), .Q (n_2498));
  ON21X1 g62735(.A (n_1601), .B (n_1685), .C (n_1864), .Q (n_2497));
  NA2X1 g62736(.A (n_2318), .B (n_2319), .Q (n_2496));
  AN22X1 g62737(.A (n_2169), .B (n_5317), .C (n_2167), .D (n_5318), .Q
       (n_2495));
  AN22X1 g62738(.A (n_2165), .B (n_5321), .C (n_2171), .D (n_5319), .Q
       (n_2494));
  ON21X1 g62739(.A (n_1601), .B (n_1681), .C (n_1862), .Q (n_2493));
  AN22X1 g62740(.A (n_2181), .B (n_4968), .C (n_2177), .D (n_4969), .Q
       (n_2492));
  AN22X1 g62741(.A (n_2179), .B (n_5001), .C (n_2177), .D (n_5000), .Q
       (n_2491));
  AN22X1 g62742(.A (n_2181), .B (n_4999), .C (n_2195), .D (n_5004), .Q
       (n_2490));
  AO22X1 g62743(.A (n_2191), .B (n_4944), .C (n_2183), .D (n_4940), .Q
       (n_2489));
  AO22X1 g62744(.A (n_2193), .B (n_4941), .C (n_2195), .D (n_4942), .Q
       (n_2488));
  AN22X1 g62745(.A (n_2196), .B (n_4974), .C (n_2195), .D (n_4973), .Q
       (n_2487));
  AN22X1 g62746(.A (n_2191), .B (n_4975), .C (n_2183), .D (n_4971), .Q
       (n_2486));
  AN22X1 g62747(.A (n_2193), .B (n_4972), .C (n_2179), .D (n_4970), .Q
       (n_2485));
  AN22X1 g62748(.A (n_2193), .B (n_5003), .C (n_2196), .D (n_5005), .Q
       (n_2484));
  AN22X1 g62749(.A (n_2191), .B (n_5006), .C (n_2183), .D (n_5002), .Q
       (n_2483));
  AN22X1 g62750(.A (n_2173), .B (n_4579), .C (n_2169), .D (n_4573), .Q
       (n_2482));
  AN22X1 g62751(.A (n_2200), .B (n_4990), .C (n_2153), .D (n_4992), .Q
       (n_2481));
  AN22X1 g62752(.A (n_2176), .B (n_5506), .C (n_1813), .D (n_5510), .Q
       (n_2480));
  AN22X1 g62753(.A (n_2176), .B (n_4576), .C (n_1813), .D (n_4580), .Q
       (n_2479));
  AN22X1 g62754(.A (n_2176), .B (n_5289), .C (n_1813), .D (n_5293), .Q
       (n_2478));
  ON21X1 g62755(.A (n_1601), .B (n_1665), .C (n_1860), .Q (n_2477));
  AN22X1 g62756(.A (n_2154), .B (n_4936), .C (n_2156), .D (n_4935), .Q
       (n_2476));
  AN22X1 g62757(.A (n_2150), .B (n_4932), .C (n_2152), .D (n_4931), .Q
       (n_2475));
  NO2X1 g62758(.A (n_2334), .B (n_2335), .Q (n_2474));
  AN21X1 g62759(.A (n_2154), .B (n_4998), .C (n_2333), .Q (n_2473));
  AN22X1 g62760(.A (n_2150), .B (n_4994), .C (n_2152), .D (n_4993), .Q
       (n_2472));
  ON22X1 g62761(.A (n_2203), .B (n_1708), .C (n_2199), .D (n_1680), .Q
       (n_2471));
  AN22X1 g62762(.A (n_1595), .B (n_4894), .C (n_2188), .D (n_4891), .Q
       (n_2470));
  AN22X1 g62763(.A (n_2185), .B (n_4893), .C (n_2187), .D (n_4892), .Q
       (n_2469));
  AN22X1 g62764(.A (n_2179), .B (n_4908), .C (n_2177), .D (n_4907), .Q
       (n_2468));
  AN22X1 g62765(.A (n_2191), .B (n_4913), .C (n_2183), .D (n_4909), .Q
       (n_2467));
  AN22X1 g62766(.A (n_2196), .B (n_4912), .C (n_2181), .D (n_4906), .Q
       (n_2466));
  AN22X1 g62767(.A (n_2193), .B (n_4910), .C (n_2195), .D (n_4911), .Q
       (n_2465));
  AN21X1 g62768(.A (n_2154), .B (n_4905), .C (n_2328), .Q (n_2464));
  AN22X1 g62769(.A (n_2200), .B (n_4897), .C (n_2153), .D (n_4899), .Q
       (n_2463));
  AN21X1 g62771(.A (n_2176), .B (n_5165), .C (n_1905), .Q (n_2462));
  AN22X1 g62772(.A (n_2176), .B (n_5041), .C (n_1813), .D (n_5045), .Q
       (n_2461));
  ON21X1 g62773(.A (n_1601), .B (n_1711), .C (n_1827), .Q (n_2460));
  ON21X1 g62774(.A (n_1601), .B (n_1682), .C (n_1835), .Q (n_2459));
  AN22X1 g62775(.A (n_2169), .B (n_4945), .C (n_2167), .D (n_4946), .Q
       (n_2458));
  AN22X1 g62776(.A (n_2165), .B (n_4949), .C (n_2171), .D (n_4947), .Q
       (n_2457));
  AN22X1 g62777(.A (n_2173), .B (n_4982), .C (n_2169), .D (n_4976), .Q
       (n_2456));
  AN22X1 g62778(.A (n_2165), .B (n_4980), .C (n_1600), .D (n_4981), .Q
       (n_2455));
  AN22X1 g62779(.A (n_2173), .B (n_5013), .C (n_1600), .D (n_5012), .Q
       (n_2454));
  AN22X1 g62780(.A (n_2169), .B (n_5007), .C (n_2171), .D (n_5009), .Q
       (n_2453));
  AN22X1 g62781(.A (n_2165), .B (n_5011), .C (n_2167), .D (n_5008), .Q
       (n_2452));
  NO2X1 g62782(.A (n_2309), .B (n_2310), .Q (n_2451));
  AN21X1 g62783(.A (n_2154), .B (n_4874), .C (n_2308), .Q (n_2450));
  NO2X1 g62784(.A (n_2305), .B (n_2306), .Q (n_2449));
  NO2X1 g62785(.A (n_2312), .B (n_2307), .Q (n_2448));
  AN21X1 g62786(.A (n_2188), .B (n_4860), .C (n_2317), .Q (n_2447));
  NO2X1 g62787(.A (n_2315), .B (n_2316), .Q (n_2446));
  NO2X1 g62788(.A (n_2313), .B (n_2314), .Q (n_2445));
  NA2X1 g62789(.A (n_2301), .B (n_2302), .Q (n_2444));
  AO22X1 g62790(.A (n_2191), .B (n_4882), .C (n_2183), .D (n_4878), .Q
       (n_2443));
  AN22X1 g62791(.A (n_2181), .B (n_4875), .C (n_2177), .D (n_4876), .Q
       (n_2442));
  AN22X1 g62792(.A (n_2173), .B (n_4920), .C (n_1598), .D (n_4919), .Q
       (n_2441));
  AN22X1 g62793(.A (n_2169), .B (n_4914), .C (n_2167), .D (n_4915), .Q
       (n_2440));
  AN22X1 g62794(.A (n_2165), .B (n_4918), .C (n_2171), .D (n_4916), .Q
       (n_2439));
  AN22X1 g62795(.A (n_2193), .B (n_4879), .C (n_2195), .D (n_4880), .Q
       (n_2438));
  AN22X1 g62798(.A (n_2150), .B (n_4777), .C (n_2152), .D (n_4776), .Q
       (n_2435));
  AN22X1 g62799(.A (n_2200), .B (n_4773), .C (n_2153), .D (n_4775), .Q
       (n_2434));
  ON22X1 g62800(.A (n_1594), .B (n_1704), .C (n_2189), .D (n_1673), .Q
       (n_2433));
  AN22X1 g62801(.A (n_2185), .B (n_4769), .C (n_2187), .D (n_4768), .Q
       (n_2432));
  AN22X1 g62802(.A (n_2202), .B (n_4772), .C (n_2198), .D (n_4771), .Q
       (n_2431));
  NO2X1 g62803(.A (n_2299), .B (n_2300), .Q (n_2430));
  NO2X1 g62804(.A (n_2296), .B (n_2298), .Q (n_2429));
  NO2X1 g62805(.A (n_2295), .B (n_2297), .Q (n_2428));
  AN22X1 g62806(.A (n_2193), .B (n_4786), .C (n_2195), .D (n_4787), .Q
       (n_2427));
  NO2X1 g62807(.A (n_2292), .B (n_2293), .Q (n_2426));
  NO2X1 g62808(.A (n_2290), .B (n_2291), .Q (n_2425));
  AN22X1 g62809(.A (n_2165), .B (n_4887), .C (n_1600), .D (n_4888), .Q
       (n_2424));
  ON21X1 g62810(.A (n_1601), .B (n_1706), .C (n_1834), .Q (n_2423));
  ON21X1 g62811(.A (n_1601), .B (n_1709), .C (n_1826), .Q (n_2422));
  AN22X1 g62812(.A (n_2176), .B (n_5010), .C (n_1813), .D (n_5014), .Q
       (n_2421));
  NO2X1 g62813(.A (n_2286), .B (n_2287), .Q (n_2420));
  NO2X1 g62814(.A (n_2284), .B (n_2285), .Q (n_2419));
  NO2X1 g62815(.A (n_2282), .B (n_2283), .Q (n_2418));
  AN21X1 g62816(.A (n_2176), .B (n_4917), .C (n_1833), .Q (n_2417));
  AN22X1 g62818(.A (n_2179), .B (n_4815), .C (n_2177), .D (n_4814), .Q
       (n_2415));
  AN22X1 g62819(.A (n_2185), .B (n_4800), .C (n_2187), .D (n_4799), .Q
       (n_2414));
  AN22X1 g62820(.A (n_2147), .B (n_4801), .C (n_2188), .D (n_4798), .Q
       (n_2413));
  AN22X1 g62821(.A (n_2191), .B (n_4820), .C (n_2183), .D (n_4816), .Q
       (n_2412));
  AN22X1 g62822(.A (n_2196), .B (n_4819), .C (n_2181), .D (n_4813), .Q
       (n_2411));
  AN22X1 g62823(.A (n_2147), .B (n_4739), .C (n_2188), .D (n_4736), .Q
       (n_2410));
  AN22X1 g62824(.A (n_2185), .B (n_4738), .C (n_2187), .D (n_4737), .Q
       (n_2409));
  NO2X1 g62825(.A (n_2280), .B (n_2281), .Q (n_2408));
  AN22X1 g62826(.A (n_2191), .B (n_4758), .C (n_2183), .D (n_4754), .Q
       (n_2407));
  NO2X1 g62827(.A (n_2278), .B (n_2279), .Q (n_2406));
  AN22X1 g62828(.A (n_2193), .B (n_4817), .C (n_2195), .D (n_4818), .Q
       (n_2405));
  AN22X1 g62829(.A (n_2202), .B (n_4741), .C (n_2198), .D (n_4740), .Q
       (n_2404));
  NO2X1 g62830(.A (n_2276), .B (n_2277), .Q (n_2403));
  AN22X1 g62831(.A (n_2202), .B (n_4803), .C (n_2198), .D (n_4802), .Q
       (n_2402));
  AN22X1 g62832(.A (n_2200), .B (n_4804), .C (n_2153), .D (n_4806), .Q
       (n_2401));
  AN22X1 g62833(.A (n_2200), .B (n_4742), .C (n_2153), .D (n_4744), .Q
       (n_2400));
  AN22X1 g62835(.A (n_2171), .B (n_4823), .C (n_2167), .D (n_4822), .Q
       (n_2398));
  NO2X1 g62837(.A (n_2269), .B (n_2270), .Q (n_2396));
  NO2X1 g62838(.A (n_2267), .B (n_2268), .Q (n_2395));
  NO2X1 g62839(.A (n_2273), .B (n_2274), .Q (n_2394));
  AN22X1 g62840(.A (n_2173), .B (n_4827), .C (n_2169), .D (n_4821), .Q
       (n_2393));
  AN22X1 g62842(.A (n_2154), .B (n_4812), .C (n_2156), .D (n_4811), .Q
       (n_2391));
  AN22X1 g62843(.A (n_2150), .B (n_4808), .C (n_2152), .D (n_4807), .Q
       (n_2390));
  AN22X1 g62845(.A (n_2154), .B (n_4750), .C (n_2156), .D (n_4749), .Q
       (n_2388));
  AN22X1 g62846(.A (n_2150), .B (n_4746), .C (n_2152), .D (n_4745), .Q
       (n_2387));
  AN21X1 g62847(.A (n_2176), .B (n_4824), .C (n_1829), .Q (n_2386));
  ON21X1 g62848(.A (n_1601), .B (n_1672), .C (n_1828), .Q (n_2385));
  AND6X1 g62849(.A (n_2289), .B (n_1927), .C (n_1928), .D (n_2020), .E
       (n_1916), .F (n_1925), .Q (n_2590));
  NA2X1 g62850(.A (n_2383), .B (n_2018), .Q (n_2589));
  NA2X1 g62851(.A (n_2384), .B (n_2018), .Q (n_2588));
  NA2X1 g62852(.A (n_2383), .B (n_2019), .Q (n_2587));
  NA2X1 g62853(.A (n_2384), .B (n_2019), .Q (n_2586));
  INX1 g62854(.A (n_2384), .Q (n_2383));
  HAX1 g62855(.A (n_2010), .B (n_1700), .S (n_2384), .CO (n_2379));
  NO2I1X1 g62856(.B (n_2172), .AN (n_5164), .Q (n_2378));
  NO2I1X1 g62857(.B (n_2166), .AN (n_5228), .Q (n_2377));
  NO2I1X1 g62858(.B (n_2172), .AN (n_5226), .Q (n_2376));
  AN221X1 g62859(.A (csr_mcause[15]), .B (n_2012), .C (n_2016), .D
       (csr_mtval[15]), .E (n_2230), .Q (n_2375));
  AN221X1 g62860(.A (csr_mscratch[13]), .B (n_1970), .C (n_2014), .D
       (n_5553), .E (n_2208), .Q (n_2374));
  AN221X1 g62861(.A (csr_mscratch[14]), .B (n_1970), .C (n_2014), .D
       (n_5552), .E (n_2209), .Q (n_2373));
  AN221X1 g62863(.A (csr_mscratch[10]), .B (n_1970), .C (n_2014), .D
       (n_5557), .E (n_2137), .Q (n_2371));
  AN221X1 g62864(.A (csr_mscratch[9]), .B (n_1970), .C (n_2014), .D
       (n_5558), .E (n_2135), .Q (n_2370));
  NO2I1X1 g62865(.B (n_2158), .AN (n_5522), .Q (n_2369));
  NO2I1X1 g62866(.B (n_2158), .AN (n_5460), .Q (n_2368));
  NO2I1X1 g62868(.B (n_2158), .AN (n_5181), .Q (n_2366));
  NO2I1X1 g62869(.B (n_1594), .AN (n_5049), .Q (n_2365));
  NO2I1X1 g62870(.B (n_2163), .AN (n_5275), .Q (n_2364));
  NO2I1X1 g62871(.B (n_2158), .AN (n_5398), .Q (n_2363));
  NO2I1X1 g62874(.B (n_2158), .AN (n_5243), .Q (n_2360));
  AN221X1 g62875(.A (csr_mscratch[6]), .B (n_1970), .C (n_2014), .D
       (n_5561), .E (n_2129), .Q (n_2359));
  NO2I1X1 g62876(.B (n_2158), .AN (n_5491), .Q (n_2358));
  NO2I1X1 g62877(.B (n_2158), .AN (n_4561), .Q (n_2357));
  NO2I1X1 g62878(.B (n_2189), .AN (n_5139), .Q (n_2356));
  NO2I1X1 g62879(.B (n_2189), .AN (n_5015), .Q (n_2355));
  NO2I1X1 g62880(.B (n_1594), .AN (n_5142), .Q (n_2354));
  NO2I1X1 g62881(.B (n_1594), .AN (n_5018), .Q (n_2353));
  NA2X1 g62883(.A (n_2164), .B (n_5213), .Q (n_2351));
  NA2X1 g62884(.A (n_2164), .B (n_5151), .Q (n_2350));
  NA2X1 g62885(.A (n_2164), .B (n_5027), .Q (n_2349));
  NO2I1X1 g62886(.B (n_2157), .AN (n_5214), .Q (n_2348));
  NO2I1X1 g62887(.B (n_2155), .AN (n_5215), .Q (n_2347));
  NO2I1X1 g62888(.B (n_1597), .AN (n_5022), .Q (n_2346));
  NO2I1X1 g62889(.B (n_2158), .AN (n_5026), .Q (n_2345));
  NO2I1X1 g62891(.B (n_2158), .AN (n_5305), .Q (n_2343));
  NO2I1X1 g62893(.B (n_1597), .AN (n_4960), .Q (n_2341));
  NO2I1X1 g62894(.B (n_2158), .AN (n_4964), .Q (n_2340));
  NO2I1X1 g62896(.B (n_1597), .AN (n_4929), .Q (n_2338));
  NO2I1X1 g62897(.B (n_2158), .AN (n_4933), .Q (n_2337));
  NA2X1 g62898(.A (n_2164), .B (n_4996), .Q (n_2336));
  NO2I1X1 g62899(.B (n_2162), .AN (n_4991), .Q (n_2335));
  NO2I1X1 g62900(.B (n_2158), .AN (n_4995), .Q (n_2334));
  NO2I1X1 g62901(.B (n_2157), .AN (n_4997), .Q (n_2333));
  NO2I1X1 g62902(.B (n_2148), .AN (n_4987), .Q (n_2332));
  AN221X1 g62903(.A (csr_mscratch[5]), .B (n_1970), .C (n_2014), .D
       (n_5562), .E (n_2128), .Q (n_2331));
  NO2I1X1 g62904(.B (n_1597), .AN (n_4898), .Q (n_2330));
  NO2I1X1 g62905(.B (n_2158), .AN (n_4902), .Q (n_2329));
  NO2I1X1 g62906(.B (n_2157), .AN (n_4904), .Q (n_2328));
  NO2I1X1 g62907(.B (n_2175), .AN (n_5229), .Q (n_2327));
  NO2I1X1 g62908(.B (n_2174), .AN (n_5230), .Q (n_2326));
  NO2I1X1 g62909(.B (n_2168), .AN (n_5225), .Q (n_2325));
  NO2I1X1 g62910(.B (n_2170), .AN (n_5224), .Q (n_2324));
  NO2X1 g62911(.A (n_6067), .B (n_1841), .Q (n_2382));
  OR2X1 g62912(.A (n_6064), .B (n_1841), .Q (n_2381));
  ON21X1 g62913(.A (n_5573), .B (n_1854), .C (n_1906), .Q (n_2380));
  INX1 g62914(.A (n_2322), .Q (n_2323));
  NO2I1X1 g62915(.B (n_2174), .AN (n_5168), .Q (n_2320));
  NA2X1 g62916(.A (n_1598), .B (n_5353), .Q (n_2319));
  NA2X1 g62917(.A (n_2169), .B (n_5348), .Q (n_2318));
  NO2I1X1 g62918(.B (n_2148), .AN (n_4863), .Q (n_2317));
  NO2I1X1 g62919(.B (n_2186), .AN (n_4861), .Q (n_2316));
  NO2I1X1 g62920(.B (n_2184), .AN (n_4862), .Q (n_2315));
  NO2I1X1 g62921(.B (n_2199), .AN (n_4864), .Q (n_2314));
  NO2I1X1 g62922(.B (n_2203), .AN (n_4865), .Q (n_2313));
  NO2I1X1 g62923(.B (n_2201), .AN (n_4866), .Q (n_2312));
  NA2X1 g62924(.A (n_2164), .B (n_4872), .Q (n_2311));
  NO2I1X1 g62925(.B (n_2162), .AN (n_4867), .Q (n_2310));
  NO2I1X1 g62926(.B (n_2158), .AN (n_4871), .Q (n_2309));
  NO2I1X1 g62927(.B (n_2157), .AN (n_4873), .Q (n_2308));
  NO2I1X1 g62928(.B (n_1573), .AN (n_4868), .Q (n_2307));
  NO2I1X1 g62929(.B (n_2151), .AN (n_4869), .Q (n_2306));
  NO2I1X1 g62930(.B (n_2149), .AN (n_4870), .Q (n_2305));
  AN222X1 g62931(.A (n_3263), .B (n_2017), .C (n_4549), .D (n_5723), .E
       (n_1936), .F (csr_mtvec[7]), .Q (n_2304));
  NA2X1 g62933(.A (n_2179), .B (n_4877), .Q (n_2302));
  NA2X1 g62934(.A (n_2196), .B (n_4881), .Q (n_2301));
  NO2I1X1 g62935(.B (n_2178), .AN (n_4783), .Q (n_2300));
  NO2I1X1 g62936(.B (n_2180), .AN (n_4784), .Q (n_2299));
  NO2I1X1 g62937(.B (n_1575), .AN (n_4785), .Q (n_2298));
  NO2I1X1 g62938(.B (n_2182), .AN (n_4782), .Q (n_2297));
  NO2I1X1 g62939(.B (n_2190), .AN (n_4789), .Q (n_2296));
  NO2I1X1 g62940(.B (n_2197), .AN (n_4788), .Q (n_2295));
  NO2I1X1 g62941(.B (n_1601), .AN (n_4886), .Q (n_2294));
  NO2I1X1 g62942(.B (n_2168), .AN (n_4884), .Q (n_2293));
  NO2I1X1 g62943(.B (n_2172), .AN (n_4885), .Q (n_2292));
  NO2I1X1 g62944(.B (n_2170), .AN (n_4883), .Q (n_2291));
  NO2I1X1 g62945(.B (n_2174), .AN (n_4889), .Q (n_2290));
  AND6X1 g62946(.A (n_2086), .B (n_1919), .C (n_1918), .D (n_2021), .E
       (n_1929), .F (n_1920), .Q (n_2289));
  ON21X1 g62947(.A (n_2085), .B (n_6071), .C (n_121), .Q (n_6501));
  NO2I1X1 g62948(.B (n_1601), .AN (n_4793), .Q (n_2288));
  NO2I1X1 g62949(.B (n_2175), .AN (n_4795), .Q (n_2287));
  NO2I1X1 g62950(.B (n_2174), .AN (n_4796), .Q (n_2286));
  NO2I1X1 g62951(.B (n_2168), .AN (n_4791), .Q (n_2285));
  NO2I1X1 g62952(.B (n_2170), .AN (n_4790), .Q (n_2284));
  NO2I1X1 g62953(.B (n_2172), .AN (n_4792), .Q (n_2283));
  NO2I1X1 g62954(.B (n_2166), .AN (n_4794), .Q (n_2282));
  NO2I1X1 g62955(.B (n_2178), .AN (n_4752), .Q (n_2281));
  NO2I1X1 g62956(.B (n_2180), .AN (n_4753), .Q (n_2280));
  NO2I1X1 g62957(.B (n_2182), .AN (n_4751), .Q (n_2279));
  NO2I1X1 g62958(.B (n_2197), .AN (n_4757), .Q (n_2278));
  NO2I1X1 g62959(.B (n_2194), .AN (n_4756), .Q (n_2277));
  NO2I1X1 g62960(.B (n_2192), .AN (n_4755), .Q (n_2276));
  AN222X1 g62961(.A (n_2017), .B (n_3264), .C (csr_mscratch[3]), .D
       (n_1970), .E (csr_mcycle[35]), .F (n_1937), .Q (n_2275));
  NO2I1X1 g62962(.B (n_2175), .AN (n_4826), .Q (n_2274));
  NO2I1X1 g62963(.B (n_2166), .AN (n_4825), .Q (n_2273));
  NO2I1X1 g62966(.B (n_2168), .AN (n_4760), .Q (n_2270));
  NO2I1X1 g62967(.B (n_2170), .AN (n_4759), .Q (n_2269));
  NO2I1X1 g62968(.B (n_2172), .AN (n_4761), .Q (n_2268));
  NO2I1X1 g62969(.B (n_2166), .AN (n_4763), .Q (n_2267));
  NO2X1 g62972(.A (n_2205), .B (\instruction[7]_39562 ), .Q (n_2322));
  NA2X1 g62973(.A (n_2204), .B (\instruction[7]_39562 ), .Q (n_2321));
  INX1 g62974(.A (n_6461), .Q (n_2264));
  INX1 g62975(.A (n_2263), .Q (n_2262));
  AN22X1 g62976(.A (n_2014), .B (n_5550), .C (n_2012), .D
       (csr_mcause[16]), .Q (n_2261));
  AN22X1 g62977(.A (n_2017), .B (n_3270), .C (n_1970), .D
       (csr_mscratch[21]), .Q (n_2260));
  AN22X1 g62978(.A (n_2017), .B (n_3268), .C (n_1970), .D
       (csr_mscratch[19]), .Q (n_2259));
  AN22X1 g62979(.A (n_2017), .B (n_3274), .C (n_1970), .D
       (csr_mscratch[25]), .Q (n_2258));
  AN22X1 g62980(.A (n_2017), .B (n_3271), .C (n_1970), .D
       (csr_mscratch[22]), .Q (n_2257));
  AN221X1 g62981(.A (csr_minstret[30]), .B (n_6625), .C (n_1938), .D
       (csr_minstret[62]), .E (n_2107), .Q (n_2256));
  AN221X1 g62982(.A (csr_mcycle[15]), .B (n_6624), .C (n_1937), .D
       (csr_mcycle[47]), .E (n_2102), .Q (n_2255));
  AN221X1 g62983(.A (csr_mcycle[13]), .B (n_6624), .C (n_1937), .D
       (csr_mcycle[45]), .E (n_2103), .Q (n_2254));
  AN221X1 g62984(.A (csr_mcycle[14]), .B (n_6624), .C (n_1937), .D
       (csr_mcycle[46]), .E (n_2104), .Q (n_2253));
  AN221X1 g62985(.A (csr_minstret[11]), .B (n_6625), .C (n_1938), .D
       (csr_minstret[43]), .E (n_2048), .Q (n_2252));
  AN221X1 g62986(.A (csr_mcycle[10]), .B (n_6624), .C (n_1937), .D
       (csr_mcycle[42]), .E (n_2056), .Q (n_2251));
  AN221X1 g62987(.A (csr_mcycle[9]), .B (n_6624), .C (n_1937), .D
       (csr_mcycle[41]), .E (n_2052), .Q (n_2250));
  AN221X1 g62988(.A (csr_mcycle[6]), .B (n_6624), .C (n_1937), .D
       (csr_mcycle[38]), .E (n_2045), .Q (n_2249));
  AN221X1 g62989(.A (csr_mcycle[5]), .B (n_6624), .C (csr_mcycle[37]),
       .D (n_1937), .E (n_2042), .Q (n_2248));
  AN22X1 g62990(.A (n_1942), .B (n_6343), .C (n_2016), .D
       (csr_mtval[30]), .Q (n_2247));
  AN22X1 g62991(.A (n_2014), .B (n_5544), .C (n_2012), .D
       (csr_mcause[22]), .Q (n_2246));
  AN22X1 g62992(.A (n_2014), .B (n_5543), .C (n_2012), .D
       (csr_mcause[31]), .Q (n_2245));
  AN22X1 g62993(.A (n_2014), .B (n_5546), .C (n_2012), .D
       (csr_mcause[20]), .Q (n_2244));
  AN22X1 g62994(.A (n_2014), .B (n_5554), .C (n_2012), .D
       (csr_mcause[30]), .Q (n_2243));
  AN22X1 g62995(.A (n_2014), .B (n_5565), .C (n_2012), .D
       (csr_mcause[29]), .Q (n_2242));
  AN22X1 g62996(.A (n_2014), .B (n_5567), .C (n_2012), .D
       (csr_mcause[28]), .Q (n_2241));
  AN22X1 g62997(.A (n_2014), .B (n_5568), .C (n_2012), .D
       (csr_mcause[27]), .Q (n_2240));
  AN22X1 g62998(.A (n_2014), .B (n_5569), .C (n_2012), .D
       (csr_mcause[26]), .Q (n_2239));
  AN22X1 g62999(.A (n_2014), .B (n_5570), .C (n_2012), .D
       (csr_mcause[25]), .Q (n_2238));
  AN22X1 g63000(.A (n_2014), .B (n_5571), .C (n_2012), .D
       (csr_mcause[24]), .Q (n_2237));
  AN22X1 g63001(.A (n_2014), .B (n_5572), .C (n_2012), .D
       (csr_mcause[23]), .Q (n_2236));
  AN22X1 g63002(.A (n_2014), .B (n_5545), .C (n_2012), .D
       (csr_mcause[21]), .Q (n_2235));
  AN22X1 g63003(.A (n_2014), .B (n_5547), .C (n_2012), .D
       (csr_mcause[19]), .Q (n_2234));
  AN22X1 g63004(.A (n_2014), .B (n_5548), .C (n_2012), .D
       (csr_mcause[18]), .Q (n_2233));
  AN22X1 g63005(.A (n_2014), .B (n_5549), .C (n_2012), .D
       (csr_mcause[17]), .Q (n_2232));
  AN22X1 g63006(.A (n_2017), .B (n_3272), .C (n_1970), .D
       (csr_mscratch[23]), .Q (n_2231));
  AO22X1 g63007(.A (n_1970), .B (csr_mscratch[15]), .C (n_2014), .D
       (n_5551), .Q (n_2230));
  AN222X1 g63008(.A (csr_utime[28]), .B (n_1837), .C (csr_utime[60]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[28]), .Q (n_2229));
  AN222X1 g63009(.A (csr_utime[31]), .B (n_1837), .C (csr_utime[63]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[31]), .Q (n_2228));
  AN222X1 g63010(.A (csr_utime[29]), .B (n_1837), .C (csr_utime[61]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[29]), .Q (n_2227));
  AN222X1 g63011(.A (csr_utime[27]), .B (n_1837), .C (csr_utime[59]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[27]), .Q (n_2226));
  AN222X1 g63012(.A (csr_utime[26]), .B (n_1837), .C (csr_utime[58]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[26]), .Q (n_2225));
  AN222X1 g63013(.A (csr_utime[25]), .B (n_1837), .C (csr_utime[57]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[25]), .Q (n_2224));
  AN222X1 g63014(.A (csr_utime[24]), .B (n_1837), .C (csr_utime[56]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[24]), .Q (n_2223));
  AN222X1 g63015(.A (csr_utime[23]), .B (n_1837), .C (csr_utime[55]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[23]), .Q (n_2222));
  AN222X1 g63016(.A (csr_utime[22]), .B (n_1837), .C (csr_utime[54]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[22]), .Q (n_2221));
  AN222X1 g63017(.A (csr_utime[21]), .B (n_1837), .C (csr_utime[53]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[21]), .Q (n_2220));
  AN222X1 g63018(.A (csr_utime[19]), .B (n_1837), .C (csr_utime[51]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[19]), .Q (n_2219));
  AN222X1 g63019(.A (csr_utime[18]), .B (n_1837), .C (csr_utime[50]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[18]), .Q (n_2218));
  AN222X1 g63020(.A (csr_utime[20]), .B (n_1837), .C (csr_utime[52]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[20]), .Q (n_2217));
  AN222X1 g63021(.A (csr_utime[17]), .B (n_1837), .C (csr_utime[49]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[17]), .Q (n_2216));
  AN222X1 g63022(.A (csr_utime[16]), .B (n_1837), .C (csr_utime[48]),
       .D (n_1836), .E (n_2016), .F (csr_mtval[16]), .Q (n_2215));
  AN22X1 g63023(.A (n_2017), .B (n_3280), .C (n_1970), .D
       (csr_mscratch[31]), .Q (n_2214));
  AN22X1 g63024(.A (n_2017), .B (n_3279), .C (n_1970), .D
       (csr_mscratch[30]), .Q (n_2213));
  AN22X1 g63025(.A (n_2017), .B (n_3278), .C (n_1970), .D
       (csr_mscratch[29]), .Q (n_2212));
  AN22X1 g63026(.A (n_2017), .B (n_3277), .C (n_1970), .D
       (csr_mscratch[28]), .Q (n_2211));
  AN22X1 g63027(.A (n_2017), .B (n_3276), .C (n_1970), .D
       (csr_mscratch[27]), .Q (n_2210));
  AO22X1 g63028(.A (n_2012), .B (csr_mcause[14]), .C (n_2016), .D
       (csr_mtval[14]), .Q (n_2209));
  AO22X1 g63029(.A (n_2012), .B (csr_mcause[13]), .C (n_2016), .D
       (csr_mtval[13]), .Q (n_2208));
  AN22X1 g63030(.A (n_2017), .B (n_3275), .C (n_1970), .D
       (csr_mscratch[26]), .Q (n_2207));
  AN22X1 g63031(.A (n_2017), .B (n_3273), .C (n_1970), .D
       (csr_mscratch[24]), .Q (n_2206));
  NA2X1 g63032(.A (n_5573), .B (n_5604), .Q (n_6064));
  NA2X1 g63033(.A (n_5573), .B (n_2117), .Q (n_6065));
  NA2X1 g63034(.A (n_204), .B (n_5604), .Q (n_6067));
  NO2X1 g63035(.A (n_5573), .B (n_5604), .Q (n_6461));
  NO2X1 g63036(.A (n_204), .B (n_1854), .Q (n_2263));
  INX1 g63037(.A (n_2204), .Q (n_2205));
  INX4 g63038(.A (n_2203), .Q (n_2202));
  INX4 g63039(.A (n_2201), .Q (n_2200));
  INX4 g63040(.A (n_2199), .Q (n_2198));
  INX4 g63041(.A (n_2197), .Q (n_2196));
  INX6 g63042(.A (n_2194), .Q (n_2195));
  INX4 g63043(.A (n_2192), .Q (n_2193));
  INX4 g63044(.A (n_2190), .Q (n_2191));
  INX4 g63045(.A (n_2189), .Q (n_2188));
  INX4 g63046(.A (n_2186), .Q (n_2187));
  INX8 g63047(.A (n_2184), .Q (n_2185));
  INX4 g63048(.A (n_1575), .Q (n_2183));
  INX4 g63049(.A (n_2182), .Q (n_2181));
  INX6 g63050(.A (n_2180), .Q (n_2179));
  INX4 g63051(.A (n_2178), .Q (n_2177));
  INX4 g63062(.A (n_1599), .Q (n_1600));
  INX6 g63066(.A (n_2174), .Q (n_2173));
  INX3 g63067(.A (n_2172), .Q (n_2171));
  INX3 g63068(.A (n_2170), .Q (n_2169));
  INX4 g63069(.A (n_2168), .Q (n_2167));
  INX3 g63070(.A (n_2166), .Q (n_2165));
  INX4 g63071(.A (n_2163), .Q (n_2164));
  INX1 g63072(.A (n_2162), .Q (n_2161));
  INX3 g63084(.A (n_1597), .Q (n_2160));
  INX3 g63090(.A (n_2157), .Q (n_2156));
  INX4 g63091(.A (n_2155), .Q (n_2154));
  INX4 g63092(.A (n_1573), .Q (n_2153));
  INX6 g63093(.A (n_2151), .Q (n_2152));
  INX4 g63094(.A (n_2149), .Q (n_2150));
  INX1 g63101(.A (n_1594), .Q (n_1595));
  INX1 g63105(.A (n_2148), .Q (n_2147));
  AN211X1 g63106(.A (n_1931), .B (n_1746), .C (n_1948), .D (n_1932), .Q
       (n_2146));
  AN22X1 g63107(.A (n_2017), .B (n_3267), .C (n_1970), .D
       (csr_mscratch[18]), .Q (n_2145));
  AN22X1 g63108(.A (n_2017), .B (n_3266), .C (n_1970), .D
       (csr_mscratch[17]), .Q (n_2144));
  AN22X1 g63109(.A (n_2017), .B (n_3265), .C (n_1970), .D
       (csr_mscratch[16]), .Q (n_2143));
  AN22X1 g63110(.A (n_2014), .B (n_5555), .C (n_2012), .D
       (csr_mcause[12]), .Q (n_2142));
  AN22X1 g63111(.A (n_1970), .B (csr_mscratch[12]), .C (n_2016), .D
       (csr_mtval[12]), .Q (n_2141));
  AN221X1 g63112(.A (csr_mcycle[0]), .B (n_6624), .C (csr_mcycle[32]),
       .D (n_1937), .E (n_2027), .Q (n_2140));
  ON21X1 g63113(.A (n_1969), .B (n_1565), .C (n_121), .Q (n_6472));
  AN22X1 g63114(.A (n_2014), .B (n_5556), .C (n_2012), .D
       (csr_mcause[11]), .Q (n_2139));
  ON221X1 g63115(.A (n_1565), .B (n_2011), .C (n_6071), .D (n_6373), .E
       (n_121), .Q (n_6500));
  AN22X1 g63116(.A (n_1942), .B (n_6322), .C (n_2016), .D
       (csr_mtval[11]), .Q (n_2138));
  AO22X1 g63117(.A (n_2012), .B (csr_mcause[10]), .C (n_2016), .D
       (csr_mtval[10]), .Q (n_2137));
  AN22X1 g63118(.A (n_2017), .B (n_3262), .C (n_1970), .D
       (csr_mscratch[11]), .Q (n_2136));
  AO22X1 g63119(.A (n_2012), .B (csr_mcause[9]), .C (n_2016), .D
       (csr_mtval[9]), .Q (n_2135));
  AN22X1 g63120(.A (n_1970), .B (csr_mscratch[8]), .C (n_2014), .D
       (n_5559), .Q (n_2134));
  AN222X1 g63121(.A (n_5723), .B (n_5542), .C (csr_utime[3]), .D
       (n_1837), .E (n_6325), .F (n_1942), .Q (n_2133));
  AN22X1 g63122(.A (n_2012), .B (csr_mcause[8]), .C (n_2016), .D
       (csr_mtval[8]), .Q (n_2132));
  AN22X1 g63123(.A (n_1970), .B (csr_mscratch[7]), .C (n_2014), .D
       (n_5560), .Q (n_2131));
  AN22X1 g63124(.A (n_2012), .B (csr_mcause[7]), .C (n_2016), .D
       (csr_mtval[7]), .Q (n_2130));
  AO22X1 g63125(.A (n_2012), .B (csr_mcause[6]), .C (n_2016), .D
       (csr_mtval[6]), .Q (n_2129));
  AO22X1 g63126(.A (n_2012), .B (csr_mcause[5]), .C (n_2016), .D
       (csr_mtval[5]), .Q (n_2128));
  AN22X1 g63127(.A (n_1970), .B (csr_mscratch[4]), .C (n_2014), .D
       (n_5563), .Q (n_2127));
  AN22X1 g63128(.A (n_2012), .B (csr_mcause[4]), .C (n_2016), .D
       (csr_mtval[4]), .Q (n_2126));
  AN22X1 g63129(.A (n_1970), .B (csr_mscratch[2]), .C (n_2014), .D
       (n_5566), .Q (n_2125));
  AN22X1 g63130(.A (n_2012), .B (csr_mcause[1]), .C (n_2016), .D
       (csr_mtval[1]), .Q (n_2124));
  AN22X1 g63131(.A (n_2012), .B (csr_mcause[2]), .C (n_2016), .D
       (csr_mtval[2]), .Q (n_2123));
  AN21X1 g63132(.A (n_6624), .B (csr_mcycle[1]), .C (n_2023), .Q
       (n_2122));
  AN221X1 g63133(.A (csr_utime[35]), .B (n_1836), .C (n_5564), .D
       (n_2014), .E (n_1953), .Q (n_2121));
  AN22X1 g63134(.A (n_2017), .B (n_3269), .C (n_1970), .D
       (csr_mscratch[20]), .Q (n_2120));
  AN22X1 g63135(.A (n_2012), .B (csr_mcause[3]), .C (n_2016), .D
       (csr_mtval[3]), .Q (n_2119));
  AN311X1 g63136(.A (n_1859), .B (n_6562), .C (n_1821), .D (n_1723), .E
       (n_1974), .Q (n_2204));
  NA2I1X4 g63137(.B (n_1589), .AN (n_2080), .Q (n_2203));
  NA2I1X4 g63138(.B (n_1591), .AN (n_2080), .Q (n_2201));
  NA2I1X4 g63139(.B (n_1945), .AN (n_2080), .Q (n_2199));
  NA2I1X4 g63140(.B (n_1568), .AN (n_2080), .Q (n_2197));
  NA2X2 g63141(.A (n_2079), .B (n_1590), .Q (n_2194));
  NA2X4 g63142(.A (n_2079), .B (n_1946), .Q (n_2192));
  NA2I1X4 g63143(.B (n_1949), .AN (n_2080), .Q (n_2190));
  NA2I1X4 g63144(.B (n_1945), .AN (n_2081), .Q (n_2189));
  NA2I1X2 g63145(.B (n_1589), .AN (n_2081), .Q (n_2186));
  NA2I1X2 g63146(.B (n_1591), .AN (n_2081), .Q (n_2184));
  NA2I1X2 g63148(.B (n_1946), .AN (n_2081), .Q (n_2182));
  NA2I1X2 g63149(.B (n_1568), .AN (n_2081), .Q (n_2180));
  NA2I1X2 g63150(.B (n_1590), .AN (n_2081), .Q (n_2178));
  NA2X4 g63151(.A (n_1949), .B (n_2078), .Q (n_1601));
  AND2X4 g63153(.A (n_2082), .B (n_1590), .Q (n_1598));
  NA2X1 g63154(.A (n_2082), .B (n_1590), .Q (n_2175));
  NA2I1X4 g63155(.B (n_1568), .AN (n_2083), .Q (n_2174));
  NA2I1X4 g63156(.B (n_1568), .AN (n_2077), .Q (n_2172));
  NA2I1X4 g63157(.B (n_1946), .AN (n_2077), .Q (n_2170));
  NA2I1X4 g63158(.B (n_1590), .AN (n_2077), .Q (n_2168));
  NA2I1X4 g63159(.B (n_1946), .AN (n_2083), .Q (n_2166));
  NA2I1X4 g63160(.B (n_1945), .AN (n_2083), .Q (n_2163));
  OR2X2 g63161(.A (n_1951), .B (n_2077), .Q (n_2162));
  OR2X4 g63162(.A (n_1951), .B (n_2077), .Q (n_1597));
  AND2X4 g63163(.A (n_1950), .B (n_2082), .Q (n_2159));
  OR2X4 g63164(.A (n_1951), .B (n_2083), .Q (n_2158));
  OR2X4 g63165(.A (n_1588), .B (n_2083), .Q (n_2157));
  OR2X2 g63166(.A (n_1947), .B (n_2083), .Q (n_2155));
  OR2X2 g63168(.A (n_1588), .B (n_2077), .Q (n_2151));
  OR2X4 g63169(.A (n_1947), .B (n_2077), .Q (n_2149));
  NA2I1X4 g63170(.B (n_2079), .AN (n_1951), .Q (n_1594));
  NA2I1X1 g63171(.B (n_1950), .AN (n_2080), .Q (n_2148));
  INX1 g63172(.A (n_2118), .Q (n_5716));
  INX1 g63173(.A (n_2117), .Q (n_5604));
  INX1 g63174(.A (n_204), .Q (n_5573));
  AN22X1 g63175(.A (n_6624), .B (csr_mcycle[21]), .C (n_1937), .D
       (csr_mcycle[53]), .Q (n_2116));
  AN22X1 g63176(.A (n_6624), .B (csr_mcycle[22]), .C (n_1937), .D
       (csr_mcycle[54]), .Q (n_2115));
  AN22X1 g63177(.A (n_6624), .B (csr_mcycle[23]), .C (n_1937), .D
       (csr_mcycle[55]), .Q (n_2114));
  AN22X1 g63178(.A (n_6624), .B (csr_mcycle[24]), .C (n_1937), .D
       (csr_mcycle[56]), .Q (n_2113));
  AN22X1 g63179(.A (n_6624), .B (csr_mcycle[25]), .C (n_1937), .D
       (csr_mcycle[57]), .Q (n_2112));
  AN22X1 g63180(.A (n_6624), .B (csr_mcycle[26]), .C (n_1937), .D
       (csr_mcycle[58]), .Q (n_2111));
  AN22X1 g63181(.A (n_6624), .B (csr_mcycle[27]), .C (n_1937), .D
       (csr_mcycle[59]), .Q (n_2110));
  AN22X1 g63182(.A (n_6624), .B (csr_mcycle[28]), .C (n_1937), .D
       (csr_mcycle[60]), .Q (n_2109));
  AN22X1 g63183(.A (n_6624), .B (csr_mcycle[29]), .C (n_1937), .D
       (csr_mcycle[61]), .Q (n_2108));
  AO22X1 g63184(.A (n_6624), .B (csr_mcycle[30]), .C (n_1937), .D
       (csr_mcycle[62]), .Q (n_2107));
  AN22X1 g63185(.A (n_6624), .B (csr_mcycle[31]), .C (n_1937), .D
       (csr_mcycle[63]), .Q (n_2106));
  AN22X1 g63186(.A (n_6624), .B (csr_mcycle[19]), .C (n_1937), .D
       (csr_mcycle[51]), .Q (n_2105));
  ON21X1 g63187(.A (n_1935), .B (n_1565), .C (n_121), .Q (n_6465));
  AO222X1 g63188(.A (csr_utime[14]), .B (n_1837), .C (csr_mtvec[14]),
       .D (n_1936), .E (csr_utime[46]), .F (n_1836), .Q (n_2104));
  AO222X1 g63189(.A (csr_utime[13]), .B (n_1837), .C (csr_mtvec[13]),
       .D (n_1936), .E (csr_utime[45]), .F (n_1836), .Q (n_2103));
  AO222X1 g63190(.A (csr_utime[15]), .B (n_1837), .C (csr_mtvec[15]),
       .D (n_1936), .E (csr_utime[47]), .F (n_1836), .Q (n_2102));
  AN22X1 g63191(.A (n_1942), .B (n_6326), .C (n_1936), .D
       (csr_mtvec[16]), .Q (n_2101));
  AN22X1 g63192(.A (n_1942), .B (n_6331), .C (n_1936), .D
       (csr_mtvec[20]), .Q (n_2100));
  AN22X1 g63193(.A (n_1942), .B (n_6330), .C (n_1936), .D
       (csr_mtvec[19]), .Q (n_2099));
  AN22X1 g63194(.A (n_1942), .B (n_6328), .C (n_1936), .D
       (csr_mtvec[18]), .Q (n_2098));
  AN22X1 g63195(.A (n_1942), .B (n_6327), .C (n_1936), .D
       (csr_mtvec[17]), .Q (n_2097));
  AN22X1 g63196(.A (n_1942), .B (n_6332), .C (n_1936), .D
       (csr_mtvec[21]), .Q (n_2096));
  AN22X1 g63197(.A (n_1942), .B (n_6337), .C (n_1936), .D
       (csr_mtvec[25]), .Q (n_2095));
  AN22X1 g63198(.A (n_1942), .B (n_6333), .C (n_1936), .D
       (csr_mtvec[22]), .Q (n_2094));
  AN22X1 g63199(.A (n_1942), .B (n_6336), .C (n_1936), .D
       (csr_mtvec[24]), .Q (n_2093));
  AN22X1 g63200(.A (n_1942), .B (n_6338), .C (n_1936), .D
       (csr_mtvec[26]), .Q (n_2092));
  AN22X1 g63201(.A (n_1942), .B (n_6344), .C (n_1936), .D
       (csr_mtvec[31]), .Q (n_2091));
  AN22X1 g63202(.A (n_1942), .B (n_6334), .C (n_1936), .D
       (csr_mtvec[23]), .Q (n_2090));
  AN22X1 g63203(.A (n_1942), .B (n_6342), .C (n_1936), .D
       (csr_mtvec[29]), .Q (n_2089));
  AN22X1 g63204(.A (n_1942), .B (n_6339), .C (n_1936), .D
       (csr_mtvec[27]), .Q (n_2088));
  AN22X1 g63205(.A (n_1942), .B (n_6340), .C (n_1936), .D
       (csr_mtvec[28]), .Q (n_2087));
  MU2X1 g63206(.S (n_1587), .IN0 (n_6151), .IN1 (n_6152), .Q (n_5696));
  MU2X1 g63207(.S (n_1587), .IN0 (n_6143), .IN1 (n_6144), .Q (n_5688));
  MU2IX1 g63208(.S (n_1587), .IN0 (n_6179), .IN1 (n_6180), .Q (n_2118));
  MU2X1 g63209(.S (n_1587), .IN0 (n_6177), .IN1 (n_6178), .Q (n_5714));
  MU2X1 g63210(.S (n_1587), .IN0 (n_6175), .IN1 (n_6176), .Q (n_5713));
  MU2X1 g63211(.S (n_1587), .IN0 (n_6169), .IN1 (n_6170), .Q (n_5710));
  MU2X1 g63212(.S (n_1587), .IN0 (n_6173), .IN1 (n_6174), .Q (n_5712));
  MU2X1 g63213(.S (n_1587), .IN0 (n_6171), .IN1 (n_6172), .Q (n_5711));
  MU2X1 g63214(.S (n_1587), .IN0 (n_6167), .IN1 (n_6168), .Q (n_5709));
  MU2X1 g63215(.S (n_1587), .IN0 (n_6159), .IN1 (n_6160), .Q (n_5705));
  MU2X1 g63216(.S (n_1587), .IN0 (n_6165), .IN1 (n_6166), .Q (n_5708));
  MU2X1 g63217(.S (n_1587), .IN0 (n_6153), .IN1 (n_6154), .Q (n_5698));
  MU2X1 g63218(.S (n_1587), .IN0 (n_6161), .IN1 (n_6162), .Q (n_5706));
  MU2X1 g63219(.S (n_1587), .IN0 (n_6163), .IN1 (n_6164), .Q (n_5707));
  MU2X1 g63220(.S (n_1587), .IN0 (n_6157), .IN1 (n_6158), .Q (n_5702));
  MU2X1 g63221(.S (n_1587), .IN0 (n_6155), .IN1 (n_6156), .Q (n_5700));
  MU2X1 g63222(.S (n_1587), .IN0 (n_6149), .IN1 (n_6150), .Q (n_5694));
  MU2X1 g63223(.S (n_1587), .IN0 (n_6133), .IN1 (n_6134), .Q (n_5720));
  MU2X1 g63224(.S (n_1587), .IN0 (n_6131), .IN1 (n_6132), .Q (n_5719));
  MU2X1 g63225(.S (n_1587), .IN0 (n_6129), .IN1 (n_6130), .Q (n_5718));
  MU2X1 g63226(.S (n_1587), .IN0 (n_6127), .IN1 (n_6128), .Q (n_5717));
  MU2X1 g63227(.S (n_1587), .IN0 (n_6145), .IN1 (n_6146), .Q (n_5690));
  MU2X1 g63228(.S (n_1587), .IN0 (n_6137), .IN1 (n_6138), .Q (n_5722));
  MU2X1 g63229(.S (n_1587), .IN0 (n_6121), .IN1 (n_6122), .Q (n_5682));
  MU2X1 g63230(.S (n_1587), .IN0 (n_6125), .IN1 (n_6126), .Q (n_5715));
  MU2X1 g63231(.S (n_1587), .IN0 (n_6123), .IN1 (n_6124), .Q (n_5704));
  MU2X1 g63232(.S (n_1587), .IN0 (n_6141), .IN1 (n_6142), .Q (n_5686));
  MU2X1 g63233(.S (n_1587), .IN0 (n_6139), .IN1 (n_6140), .Q (n_5684));
  MU2X1 g63234(.S (n_1587), .IN0 (n_6135), .IN1 (n_6136), .Q (n_5721));
  MU2X1 g63235(.S (n_1587), .IN0 (n_6147), .IN1 (n_6148), .Q (n_5692));
  MU2IX1 g63236(.S (n_1587), .IN0 (n_6183), .IN1 (n_6184), .Q (n_2117));
  INX1 g63238(.A (n_2084), .Q (n_2085));
  INX2 g63239(.A (n_2083), .Q (n_2082));
  INX3 g63241(.A (n_2080), .Q (n_2079));
  INX2 g63242(.A (n_2077), .Q (n_2078));
  INX2 g63244(.A (n_2076), .Q (alu_operation_code_39061));
  INX1 g63258(.A (n_2076), .Q (n_1592));
  AN22X1 g63264(.A (n_6625), .B (csr_minstret[9]), .C (n_1938), .D
       (csr_minstret[41]), .Q (n_2075));
  AN22X1 g63265(.A (n_6624), .B (csr_mcycle[18]), .C (n_1937), .D
       (csr_mcycle[50]), .Q (n_2074));
  AN22X1 g63266(.A (n_6624), .B (csr_mcycle[17]), .C (n_1937), .D
       (csr_mcycle[49]), .Q (n_2073));
  AN22X1 g63267(.A (n_6625), .B (csr_minstret[16]), .C (n_1938), .D
       (csr_minstret[48]), .Q (n_2072));
  AN22X1 g63268(.A (n_6625), .B (csr_minstret[31]), .C (n_1938), .D
       (csr_minstret[63]), .Q (n_2071));
  AN22X1 g63269(.A (n_6625), .B (csr_minstret[26]), .C (n_1938), .D
       (csr_minstret[58]), .Q (n_2070));
  AN22X1 g63270(.A (n_6625), .B (csr_minstret[29]), .C (n_1938), .D
       (csr_minstret[61]), .Q (n_2069));
  AN22X1 g63271(.A (n_6625), .B (csr_minstret[27]), .C (n_1938), .D
       (csr_minstret[59]), .Q (n_2068));
  AN22X1 g63272(.A (n_6625), .B (csr_minstret[25]), .C (n_1938), .D
       (csr_minstret[57]), .Q (n_2067));
  AN22X1 g63273(.A (n_6625), .B (csr_minstret[24]), .C (n_1938), .D
       (csr_minstret[56]), .Q (n_2066));
  AN22X1 g63274(.A (n_6625), .B (csr_minstret[23]), .C (n_1938), .D
       (csr_minstret[55]), .Q (n_2065));
  AN22X1 g63275(.A (n_6625), .B (csr_minstret[22]), .C (n_1938), .D
       (csr_minstret[54]), .Q (n_2064));
  AN22X1 g63276(.A (n_6625), .B (csr_minstret[19]), .C (n_1938), .D
       (csr_minstret[51]), .Q (n_2063));
  AN22X1 g63277(.A (n_6625), .B (csr_minstret[18]), .C (n_1938), .D
       (csr_minstret[50]), .Q (n_2062));
  AN22X1 g63278(.A (n_6624), .B (csr_mcycle[16]), .C (n_1937), .D
       (csr_mcycle[48]), .Q (n_2061));
  AN22X1 g63279(.A (n_6625), .B (csr_minstret[28]), .C (n_1938), .D
       (csr_minstret[60]), .Q (n_2060));
  AN22X1 g63280(.A (n_6625), .B (csr_minstret[21]), .C (n_1938), .D
       (csr_minstret[53]), .Q (n_2059));
  AN22X1 g63281(.A (n_6625), .B (csr_minstret[17]), .C (n_1938), .D
       (csr_minstret[49]), .Q (n_2058));
  AN22X1 g63282(.A (n_6625), .B (csr_minstret[20]), .C (n_1938), .D
       (csr_minstret[52]), .Q (n_2057));
  AO222X1 g63283(.A (csr_utime[10]), .B (n_1837), .C (csr_mtvec[10]),
       .D (n_1936), .E (csr_utime[42]), .F (n_1836), .Q (n_2056));
  AN22X1 g63284(.A (n_6625), .B (csr_minstret[15]), .C (n_1938), .D
       (csr_minstret[47]), .Q (n_2055));
  AN22X1 g63285(.A (n_6625), .B (csr_minstret[14]), .C (n_1938), .D
       (csr_minstret[46]), .Q (n_2054));
  AN22X1 g63286(.A (n_1937), .B (csr_mcycle[40]), .C (n_1936), .D
       (csr_mtvec[8]), .Q (n_2053));
  AO222X1 g63287(.A (csr_utime[9]), .B (n_1837), .C (csr_mtvec[9]), .D
       (n_1936), .E (csr_utime[41]), .F (n_1836), .Q (n_2052));
  AN22X1 g63288(.A (n_6625), .B (csr_minstret[13]), .C (n_1938), .D
       (csr_minstret[45]), .Q (n_2051));
  AN22X1 g63289(.A (n_6625), .B (csr_minstret[12]), .C (n_1938), .D
       (csr_minstret[44]), .Q (n_2050));
  AN22X1 g63290(.A (n_6624), .B (csr_mcycle[12]), .C (n_1937), .D
       (csr_mcycle[44]), .Q (n_2049));
  AO22X1 g63291(.A (n_6624), .B (csr_mcycle[11]), .C (n_1937), .D
       (csr_mcycle[43]), .Q (n_2048));
  AN22X1 g63292(.A (n_6625), .B (csr_minstret[10]), .C (n_1938), .D
       (csr_minstret[42]), .Q (n_2047));
  AN221X1 g63293(.A (csr_utime[62]), .B (n_1836), .C (n_1837), .D
       (csr_utime[30]), .E (n_1954), .Q (n_2046));
  AO222X1 g63294(.A (csr_utime[6]), .B (n_1837), .C (csr_mtvec[6]), .D
       (n_1936), .E (csr_utime[38]), .F (n_1836), .Q (n_2045));
  AN22X1 g63295(.A (n_6624), .B (csr_mcycle[8]), .C (n_6625), .D
       (csr_minstret[8]), .Q (n_2044));
  AN22X1 g63296(.A (n_6624), .B (csr_mcycle[20]), .C (n_1937), .D
       (csr_mcycle[52]), .Q (n_2043));
  AO222X1 g63297(.A (csr_utime[5]), .B (n_1837), .C (csr_mtvec[5]), .D
       (n_1936), .E (csr_utime[37]), .F (n_1836), .Q (n_2042));
  AN22X1 g63298(.A (n_6625), .B (csr_minstret[6]), .C (n_1938), .D
       (csr_minstret[38]), .Q (n_2041));
  AN22X1 g63299(.A (n_6625), .B (csr_minstret[7]), .C (n_1938), .D
       (csr_minstret[39]), .Q (n_2040));
  AN22X1 g63300(.A (n_6624), .B (csr_mcycle[7]), .C (n_1937), .D
       (csr_mcycle[39]), .Q (n_2039));
  AN22X1 g63301(.A (n_6624), .B (csr_mcycle[4]), .C (n_1936), .D
       (csr_mtvec[4]), .Q (n_2038));
  AN221X1 g63302(.A (csr_utime[44]), .B (n_1836), .C (n_1837), .D
       (csr_utime[12]), .E (n_5723), .Q (n_2037));
  AN22X1 g63303(.A (n_6624), .B (csr_mcycle[2]), .C (n_1936), .D
       (csr_mtvec[2]), .Q (n_2036));
  AN221X1 g63304(.A (csr_utime[43]), .B (n_1836), .C (n_1837), .D
       (csr_utime[11]), .E (n_5723), .Q (n_2035));
  AN222X1 g63305(.A (csr_utime[7]), .B (n_1837), .C (csr_utime[39]), .D
       (n_1836), .E (n_1942), .F (n_6324), .Q (n_2034));
  ON21X1 g63306(.A (n_1941), .B (n_1565), .C (n_121), .Q (n_6464));
  AN22X1 g63307(.A (n_6625), .B (csr_minstret[5]), .C (n_1938), .D
       (csr_minstret[37]), .Q (n_2033));
  AN22X1 g63308(.A (n_6625), .B (csr_minstret[4]), .C (n_1937), .D
       (csr_mcycle[36]), .Q (n_2032));
  AN22X1 g63309(.A (n_6624), .B (csr_mcycle[3]), .C (n_1936), .D
       (csr_mtvec[3]), .Q (n_2031));
  AN22X1 g63310(.A (n_6625), .B (csr_minstret[2]), .C (n_1937), .D
       (csr_mcycle[34]), .Q (n_2030));
  AN221X1 g63311(.A (csr_utime[40]), .B (n_1836), .C (n_1837), .D
       (csr_utime[8]), .E (n_1954), .Q (n_2029));
  AN22X1 g63312(.A (n_6625), .B (csr_minstret[3]), .C (n_1938), .D
       (csr_minstret[35]), .Q (n_2028));
  AO222X1 g63313(.A (csr_utime[0]), .B (n_1837), .C (n_6345), .D
       (n_1936), .E (csr_utime[32]), .F (n_1836), .Q (n_2027));
  AN221X1 g63314(.A (csr_utime[36]), .B (n_1836), .C (csr_utime[4]), .D
       (n_1837), .E (n_1953), .Q (n_2026));
  AN221X1 g63315(.A (csr_utime[34]), .B (n_1836), .C (csr_utime[2]), .D
       (n_1837), .E (n_1952), .Q (n_2025));
  AN22X1 g63316(.A (n_6625), .B (csr_minstret[0]), .C (n_1938), .D
       (csr_minstret[32]), .Q (n_2024));
  AO221X1 g63317(.A (csr_utime[1]), .B (n_1837), .C (n_1836), .D
       (csr_utime[33]), .E (n_1952), .Q (n_2023));
  ON211X1 g63318(.A (n_1825), .B (n_1819), .C (n_1735), .D (n_1981), .Q
       (n_2022));
  AND3X1 g63319(.A (n_1922), .B (n_1917), .C (n_1921), .Q (n_2021));
  NO3I1X1 g63320(.B (n_1982), .C (n_1914), .AN (n_1909), .Q (n_2020));
  NO3I1X1 g63321(.B (n_1980), .C (n_1911), .AN (n_1924), .Q (n_2086));
  NO2I1X1 g63322(.B (n_1974), .AN (n_1823), .Q (n_2084));
  NA2X4 g63323(.A (n_1971), .B (n_1908), .Q (n_2083));
  OR2X4 g63324(.A (n_1971), .B (n_1908), .Q (n_2081));
  OR2X4 g63325(.A (n_1971), .B (n_6787), .Q (n_2080));
  NA2X4 g63326(.A (n_1971), .B (n_6787), .Q (n_2077));
  NA2X2 g63327(.A (n_1981), .B (n_6722), .Q (n_2076));
  INX1 g63328(.A (n_2019), .Q (n_2018));
  INX1 g63329(.A (n_2016), .Q (n_2015));
  INX1 g63330(.A (n_2014), .Q (n_2013));
  INX1 g63331(.A (n_2012), .Q (n_2011));
  HAX1 g63332(.A (n_1736), .B (n_1699), .S (n_2019), .CO (n_2010));
  AO222X1 g63333(.A (csr_mtvec[26]), .B (n_1796), .C (n_1797), .D
       (n_6190), .E (n_5569), .F (n_211), .Q (n_2009));
  NA2X1 g63334(.A (n_1936), .B (csr_mtvec[12]), .Q (n_2008));
  NA2X1 g63335(.A (n_1936), .B (csr_mtvec[11]), .Q (n_2007));
  NA2X1 g63336(.A (n_1938), .B (csr_minstret[40]), .Q (n_2006));
  AO222X1 g63337(.A (csr_mtvec[27]), .B (n_1796), .C (n_1797), .D
       (n_6189), .E (n_5568), .F (n_211), .Q (n_2005));
  AO222X1 g63338(.A (csr_mtvec[23]), .B (n_1796), .C (n_1797), .D
       (n_6193), .E (n_5572), .F (n_211), .Q (n_2004));
  AO222X1 g63339(.A (csr_mtvec[19]), .B (n_1796), .C (n_1797), .D
       (n_6197), .E (n_5547), .F (n_211), .Q (n_2003));
  NA2X1 g63340(.A (n_1938), .B (csr_minstret[36]), .Q (n_2002));
  NA2X1 g63341(.A (n_1938), .B (csr_minstret[34]), .Q (n_2001));
  AO222X1 g63342(.A (csr_mtvec[31]), .B (n_1796), .C (n_1797), .D
       (n_6185), .E (n_5543), .F (n_211), .Q (n_2000));
  AO222X1 g63343(.A (csr_mtvec[30]), .B (n_1796), .C (n_1797), .D
       (n_6186), .E (n_5554), .F (n_211), .Q (n_1999));
  AO222X1 g63344(.A (csr_mtvec[29]), .B (n_1796), .C (n_1797), .D
       (n_6187), .E (n_5565), .F (n_211), .Q (n_1998));
  NA2X1 g63345(.A (n_1936), .B (csr_mtvec[30]), .Q (n_1997));
  AO222X1 g63346(.A (csr_mtvec[25]), .B (n_1796), .C (n_1797), .D
       (n_6191), .E (n_5570), .F (n_211), .Q (n_1996));
  AO222X1 g63347(.A (csr_mtvec[22]), .B (n_1796), .C (n_1797), .D
       (n_6194), .E (n_5544), .F (n_211), .Q (n_1995));
  AO222X1 g63348(.A (csr_mtvec[21]), .B (n_1796), .C (n_1797), .D
       (n_6195), .E (n_5545), .F (n_211), .Q (n_1994));
  AO222X1 g63349(.A (csr_mtvec[18]), .B (n_1796), .C (n_1797), .D
       (n_6198), .E (n_5548), .F (n_211), .Q (n_1993));
  AO222X1 g63350(.A (csr_mtvec[15]), .B (n_1796), .C (n_1797), .D
       (n_6201), .E (n_5551), .F (n_211), .Q (n_1992));
  AO222X1 g63351(.A (csr_mtvec[28]), .B (n_1796), .C (n_1797), .D
       (n_6188), .E (n_5567), .F (n_211), .Q (n_1991));
  NA5I3X1 g63352(.D (n_1821), .E (n_1698), .AN (branch_type), .BN
       (jal_type), .CN (n_1807), .Q (n_1990));
  AO222X1 g63353(.A (csr_mtvec[24]), .B (n_1796), .C (n_1797), .D
       (n_6192), .E (n_5571), .F (n_211), .Q (n_1989));
  AO222X1 g63354(.A (csr_mtvec[20]), .B (n_1796), .C (n_1797), .D
       (n_6196), .E (n_5546), .F (n_211), .Q (n_1988));
  AO222X1 g63355(.A (csr_mtvec[17]), .B (n_1796), .C (n_1797), .D
       (n_6199), .E (n_5549), .F (n_211), .Q (n_1987));
  NA2X1 g63356(.A (n_6181), .B (n_1934), .Q (n_1986));
  NO2X2 g63357(.A (n_1944), .B (n_1762), .Q (n_2017));
  NO2X4 g63358(.A (n_1944), .B (n_1567), .Q (n_2016));
  NO2X4 g63359(.A (n_1944), .B (n_1755), .Q (n_2014));
  AND2X4 g63360(.A (n_1943), .B (n_1754), .Q (n_2012));
  INX1 g63361(.A (n_1978), .Q (n_1979));
  INX1 g63362(.A (n_1976), .Q (n_1977));
  INX1 g63364(.A (n_1972), .Q (n_1973));
  INX1 g63365(.A (n_1970), .Q (n_1969));
  AO222X1 g63366(.A (csr_mtvec[14]), .B (n_1796), .C (n_1797), .D
       (n_6202), .E (n_5552), .F (n_211), .Q (n_1968));
  AO222X1 g63367(.A (csr_mtvec[11]), .B (n_1796), .C (n_1797), .D
       (n_6205), .E (n_5556), .F (n_211), .Q (n_1967));
  AO222X1 g63369(.A (csr_mtvec[16]), .B (n_1796), .C (n_1797), .D
       (n_6200), .E (n_5550), .F (n_211), .Q (n_1966));
  AO222X1 g63370(.A (csr_mtvec[10]), .B (n_1796), .C (n_1797), .D
       (n_6206), .E (n_5557), .F (n_211), .Q (n_1965));
  AO222X1 g63371(.A (csr_mtvec[13]), .B (n_1796), .C (n_1797), .D
       (n_6203), .E (n_5553), .F (n_211), .Q (n_1964));
  AN222X1 g63372(.A (n_6214), .B (n_1797), .C (n_5566), .D (n_211), .E
       (n_1796), .F (csr_mtvec[2]), .Q (n_1963));
  AO222X1 g63373(.A (csr_mtvec[9]), .B (n_1796), .C (n_1797), .D
       (n_6207), .E (n_5558), .F (n_211), .Q (n_1962));
  AO222X1 g63374(.A (csr_mtvec[12]), .B (n_1796), .C (n_1797), .D
       (n_6204), .E (n_5555), .F (n_211), .Q (n_1961));
  AO222X1 g63375(.A (csr_mtvec[8]), .B (n_1796), .C (n_1797), .D
       (n_6208), .E (n_5559), .F (n_211), .Q (n_1960));
  AO222X1 g63376(.A (csr_mtvec[7]), .B (n_1796), .C (n_1797), .D
       (n_6209), .E (n_5560), .F (n_211), .Q (n_1959));
  AO222X1 g63377(.A (csr_mtvec[6]), .B (n_1796), .C (n_1797), .D
       (n_6210), .E (n_5561), .F (n_211), .Q (n_1958));
  AO222X1 g63378(.A (csr_mtvec[5]), .B (n_1796), .C (n_1797), .D
       (n_6211), .E (n_5562), .F (n_211), .Q (n_1957));
  AO222X1 g63379(.A (csr_mtvec[4]), .B (n_1796), .C (n_1797), .D
       (n_6212), .E (n_5563), .F (n_211), .Q (n_1956));
  AO222X1 g63380(.A (n_1797), .B (n_6213), .C (csr_mtvec[3]), .D
       (n_1796), .E (n_5564), .F (n_211), .Q (n_1955));
  NO2X1 g63381(.A (n_1664), .B (n_1928), .Q (n_1985));
  OR2X1 g63382(.A (n_1664), .B (n_1925), .Q (n_1984));
  NO2X1 g63383(.A (n_1927), .B (n_1664), .Q (n_1983));
  NA2X1 g63384(.A (n_1930), .B (n_1926), .Q (n_1982));
  ON21X1 g63385(.A (n_1803), .B (n_1855), .C (n_1735), .Q (n_1981));
  NA2X1 g63386(.A (n_1923), .B (n_1912), .Q (n_1980));
  NO2X1 g63387(.A (n_1664), .B (n_1909), .Q (n_1978));
  NO2X1 g63388(.A (n_1929), .B (n_1664), .Q (n_1976));
  NO2X1 g63389(.A (n_1664), .B (n_1919), .Q (n_1975));
  AN211X1 g63390(.A (prev_load_request), .B (read_response), .C
       (n_6367), .D (n_1948), .Q (n_1974));
  NO2X1 g63391(.A (n_1918), .B (n_1664), .Q (n_1972));
  NO2X4 g63392(.A (n_1933), .B (n_1584), .Q (n_1971));
  AND2X4 g63393(.A (n_1943), .B (n_1584), .Q (n_1970));
  INX1 g63399(.A (n_1944), .Q (n_1943));
  INX1 g63400(.A (n_1942), .Q (n_1941));
  INX1 g63401(.A (n_1936), .Q (n_1935));
  INX1 g63402(.A (n_1587), .Q (n_1934));
  NO2I1X2 g63403(.B (n_1764), .AN (instruction[23]), .Q (n_1933));
  AND2X1 g63404(.A (n_1842), .B (n_1734), .Q (irq_fast_response[5]));
  ON221X1 g63405(.A (n_1696), .B (n_1768), .C (n_6459), .D (n_1726), .E
       (n_1832), .Q (n_1932));
  AND2X1 g63406(.A (n_1842), .B (n_1728), .Q (irq_fast_response[13]));
  NO2X1 g63407(.A (n_1856), .B (n_1816), .Q (n_6051));
  NO2X1 g63408(.A (n_1851), .B (n_1816), .Q (n_6049));
  AND2X1 g63409(.A (n_1842), .B (n_1733), .Q (irq_fast_response[4]));
  AND2X1 g63410(.A (n_1842), .B (n_1731), .Q (irq_fast_response[12]));
  AO21X1 g63411(.A (n_1825), .B (n_1689), .C (n_1819), .Q (n_1931));
  NO2X1 g63412(.A (n_1845), .B (n_1755), .Q (n_1954));
  NO3X1 g63413(.A (n_1772), .B (n_1819), .C (n_6722), .Q (n_5724));
  NO2X1 g63414(.A (n_1853), .B (n_1753), .Q (n_1953));
  NO2X1 g63415(.A (n_1853), .B (n_1567), .Q (n_1952));
  NA2X2 g63416(.A (n_1838), .B (n_1724), .Q (n_1951));
  NO2X1 g63417(.A (n_1839), .B (n_1725), .Q (n_1950));
  AND2X4 g63418(.A (n_1839), .B (n_1730), .Q (n_1949));
  NO2I1X1 g63419(.B (n_6367), .AN (n_1855), .Q (n_1948));
  NA2X4 g63420(.A (n_1838), .B (n_1730), .Q (n_1947));
  NO2X2 g63422(.A (n_1839), .B (n_1737), .Q (n_1589));
  NO2I1X4 g63423(.B (n_1838), .AN (n_1724), .Q (n_1946));
  AND2X4 g63425(.A (n_1838), .B (n_1583), .Q (n_1945));
  NA3X1 g63426(.A (n_1820), .B (n_1757), .C (instruction[26]), .Q
       (n_1944));
  NO2X1 g63427(.A (n_1845), .B (n_1752), .Q (n_5723));
  NO2X2 g63428(.A (n_1845), .B (n_1762), .Q (n_1942));
  AND2X4 g63431(.A (n_1570), .B (n_1824), .Q (n_1938));
  AND2X4 g63432(.A (n_1570), .B (n_1822), .Q (n_1937));
  AND3X4 g63433(.A (n_1844), .B (n_1730), .C (n_1738), .Q (n_1936));
  INX1 g63435(.A (n_1916), .Q (n_1915));
  INX1 g63436(.A (n_1913), .Q (n_1914));
  INX1 g63438(.A (n_1910), .Q (n_1911));
  AND2X1 g63439(.A (n_1843), .B (n_1728), .Q (irq_fast_response[9]));
  AND2X1 g63440(.A (n_1843), .B (n_1731), .Q (irq_fast_response[8]));
  AND2X1 g63441(.A (n_1843), .B (n_1734), .Q (irq_fast_response[1]));
  AND2X1 g63442(.A (n_1843), .B (n_1733), .Q (irq_fast_response[0]));
  AND2X1 g63443(.A (n_1846), .B (n_1728), .Q (irq_fast_response[15]));
  AND2X1 g63444(.A (n_1847), .B (n_1731), .Q (irq_fast_response[10]));
  AND2X1 g63445(.A (n_1846), .B (n_1733), .Q (irq_fast_response[6]));
  AND2X1 g63446(.A (n_1847), .B (n_1733), .Q (irq_fast_response[2]));
  AND2X1 g63447(.A (n_1847), .B (n_1728), .Q (irq_fast_response[11]));
  AND2X1 g63448(.A (n_1846), .B (n_1731), .Q (irq_fast_response[14]));
  AND2X1 g63449(.A (n_1850), .B (csr_mcause_code[2]), .Q
       (irq_timer_response));
  NO2X2 g63450(.A (n_1849), .B (csr_mcause_code[2]), .Q
       (irq_software_response));
  NA2X1 g63451(.A (n_6322), .B (n_3262), .Q (n_1930));
  NA2X1 g63452(.A (n_6326), .B (n_3265), .Q (n_1929));
  NA2X1 g63453(.A (n_6340), .B (n_3277), .Q (n_1928));
  NA2X1 g63454(.A (n_6328), .B (n_3267), .Q (n_1927));
  NA2X1 g63455(.A (n_6325), .B (n_3264), .Q (n_1926));
  NA2X1 g63456(.A (n_6343), .B (n_3279), .Q (n_1925));
  NA2X1 g63457(.A (n_6337), .B (n_3274), .Q (n_1924));
  NA2X1 g63458(.A (n_6334), .B (n_3272), .Q (n_1923));
  NA2X1 g63459(.A (n_6324), .B (n_3263), .Q (n_1922));
  NA2X1 g63460(.A (n_6344), .B (n_3280), .Q (n_1921));
  NA2X1 g63461(.A (n_6342), .B (n_3278), .Q (n_1920));
  NA2X1 g63462(.A (n_6338), .B (n_3275), .Q (n_1919));
  NA2X1 g63463(.A (n_6331), .B (n_3269), .Q (n_1918));
  NA2X1 g63464(.A (n_6339), .B (n_3276), .Q (n_1917));
  NA2X1 g63465(.A (n_6327), .B (n_3266), .Q (n_1916));
  NA2X1 g63466(.A (n_6332), .B (n_3270), .Q (n_1913));
  NA2X1 g63467(.A (n_6333), .B (n_3271), .Q (n_1912));
  NA2X1 g63468(.A (n_6336), .B (n_3273), .Q (n_1910));
  NA2X1 g63469(.A (n_6330), .B (n_3268), .Q (n_1909));
  INX1 g63471(.A (n_1907), .Q (n_1906));
  NO2I1X1 g63472(.B (n_1812), .AN (n_5169), .Q (n_1905));
  ON21X1 g63473(.A (n_1775), .B (n_1720), .C (n_1766), .Q (n_1904));
  ON21X1 g63474(.A (\rs1_data[26]_39276 ), .B (n_1720), .C (n_1814), .Q
       (n_1903));
  ON21X1 g63475(.A (n_1566), .B (n_1720), .C (n_1766), .Q (n_1902));
  ON21X1 g63476(.A (n_1773), .B (n_1720), .C (n_1766), .Q (n_1901));
  ON21X1 g63477(.A (n_1774), .B (n_1720), .C (n_1766), .Q (n_1900));
  ON21X1 g63478(.A (n_4466), .B (n_1720), .C (n_1814), .Q (n_1899));
  ON21X1 g63479(.A (\rs1_data[27]_39286 ), .B (n_1720), .C (n_1814), .Q
       (n_1898));
  ON21X1 g63480(.A (alu_sra_result[31]), .B (n_1720), .C (n_1814), .Q
       (n_1897));
  ON21X1 g63481(.A (\rs1_data[29]_39336 ), .B (n_1720), .C (n_1814), .Q
       (n_1896));
  ON21X1 g63482(.A (\rs1_data[28]_39296 ), .B (n_1720), .C (n_1814), .Q
       (n_1895));
  ON21X1 g63483(.A (\rs1_data[14]_39466 ), .B (n_1720), .C (n_1814), .Q
       (n_1894));
  ON21X1 g63484(.A (\rs1_data[23]_39246 ), .B (n_1720), .C (n_1814), .Q
       (n_1893));
  ON21X1 g63485(.A (\rs1_data[22]_39546 ), .B (n_1720), .C (n_1814), .Q
       (n_1892));
  ON21X1 g63486(.A (\rs1_data[15]_39476 ), .B (n_1720), .C (n_1814), .Q
       (n_1891));
  ON21X1 g63487(.A (n_4474), .B (n_1720), .C (n_1814), .Q (n_1890));
  ON21X1 g63488(.A (\rs1_data[21]_39536 ), .B (n_1720), .C (n_1814), .Q
       (n_1889));
  ON21X1 g63489(.A (n_4477), .B (n_1720), .C (n_1814), .Q (n_1888));
  ON21X1 g63490(.A (n_4478), .B (n_1720), .C (n_1814), .Q (n_1887));
  ON21X1 g63491(.A (\rs1_data[30]_39446 ), .B (n_1720), .C (n_1814), .Q
       (n_1886));
  ON21X1 g63492(.A (n_4481), .B (n_1720), .C (n_1814), .Q (n_1885));
  ON21X1 g63493(.A (\rs1_data[24]_39256 ), .B (n_1720), .C (n_1814), .Q
       (n_1884));
  ON21X1 g63494(.A (n_4476), .B (n_1720), .C (n_1814), .Q (n_1883));
  ON21X1 g63495(.A (n_4475), .B (n_1720), .C (n_1814), .Q (n_1882));
  ON21X1 g63496(.A (n_4486), .B (n_1720), .C (n_1814), .Q (n_1881));
  ON21X1 g63497(.A (n_4480), .B (n_1720), .C (n_1814), .Q (n_1880));
  ON21X1 g63498(.A (\rs1_data[7]_39386 ), .B (n_1720), .C (n_1814), .Q
       (n_1879));
  ON21X1 g63501(.A (\rs1_data[8]_39396 ), .B (n_1720), .C (n_1814), .Q
       (n_1876));
  ON21X1 g63502(.A (\rs1_data[16]_39486 ), .B (n_1720), .C (n_1814), .Q
       (n_1875));
  ON21X1 g63503(.A (n_4487), .B (n_1720), .C (n_1814), .Q (n_1874));
  ON21X1 g63504(.A (n_4461), .B (n_1720), .C (n_1814), .Q (n_1873));
  ON21X1 g63505(.A (\rs1_data[17]_39496 ), .B (n_1720), .C (n_1814), .Q
       (n_1872));
  NA2X1 g63507(.A (n_1813), .B (n_5138), .Q (n_1870));
  NO2I1X1 g63508(.B (n_1812), .AN (n_4704), .Q (n_1869));
  NA2X1 g63509(.A (n_1813), .B (n_5479), .Q (n_1868));
  NA2X1 g63510(.A (n_1813), .B (n_5541), .Q (n_1867));
  NA2X1 g63511(.A (n_1813), .B (n_4611), .Q (n_1866));
  NA2X1 g63512(.A (n_1813), .B (n_5107), .Q (n_1865));
  NA2X1 g63513(.A (n_1813), .B (n_5386), .Q (n_1864));
  NA2X1 g63514(.A (n_1813), .B (n_5417), .Q (n_1863));
  NA2X1 g63515(.A (n_1813), .B (n_4642), .Q (n_1862));
  ON21X1 g63516(.A (n_1776), .B (n_1720), .C (n_1766), .Q (n_1861));
  NA2X1 g63517(.A (n_1813), .B (n_5262), .Q (n_1860));
  NO2X1 g63518(.A (n_6453), .B (n_201), .Q (n_1859));
  NA2X1 g63519(.A (n_1813), .B (n_5231), .Q (n_1858));
  AN21X1 g63520(.A (n_1768), .B (n_6597), .C (n_1798), .Q (n_1907));
  INX1 g63523(.A (n_1849), .Q (n_1850));
  INX1 g63524(.A (n_1845), .Q (n_1844));
  INX1 g63525(.A (n_1841), .Q (n_1840));
  NA2X1 g63527(.A (n_1813), .B (n_5324), .Q (n_1835));
  NA2X1 g63528(.A (n_1813), .B (n_4952), .Q (n_1834));
  NO2I1X1 g63529(.B (n_1812), .AN (n_4921), .Q (n_1833));
  NA2X1 g63530(.A (branch_type), .B (n_1804), .Q (n_1832));
  NO2I1X1 g63532(.B (n_1816), .AN (n_1824), .Q (n_6048));
  NO2I1X1 g63534(.B (n_1816), .AN (n_1822), .Q (n_6050));
  NO2I1X1 g63535(.B (n_1812), .AN (n_4828), .Q (n_1829));
  NA2X1 g63536(.A (n_1813), .B (n_4766), .Q (n_1828));
  AND2X1 g63537(.A (n_1801), .B (n_1761), .Q (irq_fast_response[3]));
  NO2X2 g63538(.A (n_1569), .B (n_1760), .Q (irq_fast_response[7]));
  NA2X1 g63539(.A (n_1813), .B (n_5355), .Q (n_1827));
  NA2X1 g63540(.A (n_1813), .B (n_4983), .Q (n_1826));
  NA2X1 g63541(.A (n_1818), .B (n_1584), .Q (n_1856));
  NA3I1X1 g63542(.B (n_6605), .C (n_1771), .AN (n_6454), .Q (n_1855));
  NA2X1 g63543(.A (n_6458), .B (n_1799), .Q (n_1854));
  OR4X1 g63545(.A (n_1758), .B (n_1745), .C (n_1744), .D (n_1690), .Q
       (n_1853));
  NA2X1 g63546(.A (n_1818), .B (n_1754), .Q (n_1851));
  NA2X1 g63550(.A (n_1802), .B (n_1761), .Q (n_1849));
  ON311X1 g63552(.A (n_4457), .B (n_4456), .C (n_1715), .D (n_6373), .E
       (n_5607), .Q (n_1848));
  AND2X1 g63567(.A (n_1801), .B (csr_mcause_code[1]), .Q (n_1847));
  NO2I1X1 g63568(.B (n_1569), .AN (csr_mcause_code[1]), .Q (n_1846));
  NA3I1X1 g63569(.B (n_1818), .C (n_1757), .AN (n_6719), .Q (n_1845));
  NO2X1 g63570(.A (n_1800), .B (csr_mcause_code[1]), .Q (n_1843));
  NO2X1 g63572(.A (n_1569), .B (csr_mcause_code[1]), .Q (n_1842));
  NA2X1 g63573(.A (n_6459), .B (n_1799), .Q (n_1841));
  NO2X4 g63574(.A (n_1808), .B (n_6460), .Q (n_1839));
  AND3X4 g63575(.A (n_1818), .B (n_1770), .C (n_1756), .Q (n_1837));
  AND3X4 g63576(.A (n_1770), .B (n_1759), .C (n_1756), .Q (n_1836));
  INX1 g63578(.A (n_201), .Q (n_6367));
  INX1 g63579(.A (n_1813), .Q (n_1812));
  NA2X1 g63580(.A (n_1774), .B (n_1767), .Q (n_1811));
  NA2X1 g63582(.A (n_1566), .B (n_1767), .Q (n_1809));
  NO2X2 g63583(.A (n_1750), .B (n_1690), .Q (n_1808));
  NO2I1X1 g63584(.B (n_6602), .AN (n_1763), .Q (n_1807));
  AO21X1 g63585(.A (jalr_type), .B (n_6459), .C (jal_type), .Q
       (n_1806));
  NA2X1 g63586(.A (n_3285), .B (n_121), .Q (n_6462));
  NA2X1 g63587(.A (n_1776), .B (n_1767), .Q (n_1805));
  NA2X1 g63588(.A (n_6597), .B (n_6605), .Q (n_1804));
  NA3I1X1 g63589(.B (n_6597), .C (n_1689), .AN (n_6457), .Q (n_1803));
  NO3X4 g63590(.A (n_1725), .B (n_1582), .C (instruction[24]), .Q
       (n_6460));
  NO2I1X1 g63591(.B (n_6456), .AN (n_6722), .Q (n_1825));
  AND2X1 g63592(.A (n_1754), .B (n_1759), .Q (n_1824));
  NA3I1X1 g63593(.B (n_1768), .C (store_type), .AN
       (store_commit_cycle), .Q (n_1823));
  AND2X1 g63594(.A (n_1759), .B (n_1584), .Q (n_1822));
  NO3I1X1 g63595(.B (n_1735), .C (n_1746), .AN (n_6561), .Q (n_1821));
  NO3X1 g63596(.A (n_1741), .B (n_6719), .C (instruction[24]), .Q
       (n_1820));
  OR3X1 g63597(.A (n_1758), .B (n_1743), .C (n_6719), .Q (n_1819));
  NO2X2 g63598(.A (n_1758), .B (instruction[24]), .Q (n_1818));
  NA2X2 g63600(.A (n_1757), .B (n_6719), .Q (n_1816));
  NO5I3X1 g63601(.D (instruction[2]), .E (instruction[3]), .AN
       (n_1763), .BN (n_6718), .CN (instruction[0]), .Q (n_201));
  NO2X1 g63603(.A (n_1765), .B (n_6454), .Q (n_1814));
  AND2X4 g63604(.A (n_1756), .B (n_1690), .Q (n_1813));
  INX1 g63605(.A (n_1801), .Q (n_1800));
  INX1 g63606(.A (n_1798), .Q (n_1799));
  INX1 g63607(.A (n_1585), .Q (n_6502));
  AND2X1 g63613(.A (n_121), .B (irq_fast[10]), .Q (n_1795));
  AND2X1 g63614(.A (n_121), .B (irq_fast[8]), .Q (n_1794));
  AND2X1 g63615(.A (n_121), .B (irq_fast[2]), .Q (n_1793));
  AND2X1 g63616(.A (n_121), .B (irq_fast[11]), .Q (n_1792));
  AND2X1 g63617(.A (n_121), .B (irq_fast[0]), .Q (n_1791));
  AND2X1 g63618(.A (n_121), .B (irq_software), .Q (n_1790));
  AND2X1 g63619(.A (n_121), .B (irq_fast[14]), .Q (n_1789));
  AND2X1 g63620(.A (n_121), .B (irq_fast[13]), .Q (n_1788));
  AND2X1 g63621(.A (n_121), .B (irq_fast[15]), .Q (n_1787));
  AND2X1 g63622(.A (n_121), .B (irq_fast[4]), .Q (n_1786));
  AND2X1 g63623(.A (n_121), .B (irq_fast[7]), .Q (n_1785));
  AND2X1 g63624(.A (n_121), .B (irq_fast[6]), .Q (n_1784));
  AND2X1 g63625(.A (n_121), .B (irq_fast[12]), .Q (n_1783));
  AND2X1 g63626(.A (n_121), .B (irq_timer), .Q (n_1782));
  AND2X1 g63627(.A (n_121), .B (irq_external), .Q (n_1781));
  AND2X1 g63628(.A (n_121), .B (irq_fast[1]), .Q (n_1780));
  AND2X1 g63629(.A (n_121), .B (irq_fast[3]), .Q (n_1779));
  AND2X1 g63630(.A (n_121), .B (irq_fast[5]), .Q (n_1778));
  AND2X1 g63631(.A (n_121), .B (irq_fast[9]), .Q (n_1777));
  NO2X1 g63632(.A (n_6373), .B (csr_mcause_code[4]), .Q (n_1802));
  NO3I1X1 g63633(.B (n_6373), .C (csr_mcause_code[2]), .AN
       (csr_mcause_code[4]), .Q (n_1801));
  NA2X1 g63635(.A (n_1688), .B (n_121), .Q (n_1798));
  NO2X1 g63636(.A (n_6373), .B (n_1739), .Q (n_1797));
  NO2X1 g63637(.A (n_6373), .B (n_1740), .Q (n_1796));
  NO2X2 g63638(.A (n_1688), .B (n_1748), .Q (n_1585));
  INX1 g63639(.A (n_6455), .Q (n_1771));
  INX1 g63641(.A (n_1766), .Q (n_1765));
  MU2X2 g63642(.S (\instruction[14]_40077 ), .IN0 (n_6628), .IN1
       (n_6011), .Q (n_1776));
  MU2X2 g63643(.S (\instruction[14]_40077 ), .IN0 (n_6627), .IN1
       (n_6717), .Q (n_1775));
  MU2IX1 g63644(.S (n_1687), .IN0 (n_1703), .IN1 (n_191), .Q (n_1774));
  MU2IX1 g63645(.S (n_1687), .IN0 (n_1702), .IN1 (n_203), .Q (n_1773));
  NO2X1 g63647(.A (jalr_type), .B (jal_type), .Q (n_6562));
  NA3I1X1 g63648(.B (system_type), .C (n_6459), .AN (n_6606), .Q
       (n_1772));
  NO2X1 g63651(.A (n_1743), .B (n_1745), .Q (n_1770));
  AND2X1 g63652(.A (n_5606), .B (\instruction[14]_40077 ), .Q (n_6456));
  AND2X1 g63653(.A (n_5606), .B (n_1687), .Q (n_6458));
  AO21X1 g63654(.A (\instruction[8]_40015 ), .B (\instruction[7]_39562
       ), .C (n_1736), .Q (n_1769));
  NA2X1 g63655(.A (n_1727), .B (n_1687), .Q (n_6597));
  NO2X1 g63656(.A (n_1719), .B (\instruction[14]_40077 ), .Q (n_1768));
  OR2X1 g63657(.A (n_5606), .B (n_1727), .Q (n_1767));
  NO2X1 g63658(.A (n_1727), .B (n_5605), .Q (n_1766));
  INX1 g63659(.A (n_1760), .Q (n_1761));
  INX1 g63660(.A (n_1756), .Q (n_1755));
  INX1 g63661(.A (n_1754), .Q (n_1753));
  INX1 g63662(.A (n_1584), .Q (n_1752));
  BUX4 g63665(.A (n_1750), .Q (n_1584));
  INX1 g63668(.A (n_121), .Q (n_1748));
  NO2X4 g63671(.A (n_1725), .B (instruction[22]), .Q (n_1764));
  NO3X1 g63672(.A (\instruction[5]_40139 ), .B (instruction[4]), .C
       (instruction[6]), .Q (n_1763));
  NA2X1 g63673(.A (n_1738), .B (n_1724), .Q (n_1762));
  NA2X1 g63674(.A (n_1734), .B (csr_mcause_code[1]), .Q (n_1760));
  NO3X1 g63675(.A (n_1716), .B (instruction[25]), .C (instruction[24]),
       .Q (n_1759));
  NA2X1 g63676(.A (n_1719), .B (n_1687), .Q (n_6605));
  OR2X2 g63677(.A (n_1741), .B (instruction[26]), .Q (n_1758));
  NO2X1 g63678(.A (n_1744), .B (n_6722), .Q (n_1757));
  NO2X1 g63679(.A (n_1720), .B (n_1687), .Q (n_6454));
  NO2X2 g63680(.A (n_1729), .B (n_1582), .Q (n_1756));
  NO2X1 g63681(.A (n_1737), .B (n_1582), .Q (n_1754));
  NO2X4 g63682(.A (n_1725), .B (n_1582), .Q (n_1750));
  NA3I1X1 g63683(.B (n_1742), .C (n_4457), .AN (n_4456), .Q (n_6373));
  AND3X1 g63684(.A (n_1742), .B (n_1697), .C (n_4456), .Q (n_211));
  NO2X4 g63685(.A (reset_reg), .B (reset), .Q (n_121));
  INX1 g63686(.A (n_1739), .Q (n_1740));
  INX1 g63688(.A (n_1729), .Q (n_1730));
  INX1 g63692(.A (jalr_type), .Q (n_1726));
  INX1 g63693(.A (n_1725), .Q (n_1724));
  INX1 g63694(.A (n_1723), .Q (n_6238));
  INX1 g63695(.A (n_1720), .Q (n_1719));
  NA2X1 g63696(.A (n_6010), .B (n_1686), .Q (n_1718));
  NA2X1 g63698(.A (n_6014), .B (n_1686), .Q (n_1717));
  NA2I1X1 g63706(.B (instruction[27]), .AN (instruction[26]), .Q
       (n_1716));
  NA2I1X1 g63716(.B (current_state[0]), .AN (current_state[1]), .Q
       (n_1715));
  NO2X1 g63717(.A (n_6598), .B (n_6599), .Q (n_1746));
  NA2X1 g63718(.A (n_6722), .B (n_6719), .Q (n_1745));
  NA2X1 g63719(.A (instruction[28]), .B (instruction[29]), .Q (n_1744));
  OR2X1 g63720(.A (instruction[28]), .B (instruction[29]), .Q (n_1743));
  NO2X1 g63721(.A (current_state[0]), .B (current_state[1]), .Q
       (n_1742));
  OR2X2 g63722(.A (instruction[27]), .B (instruction[25]), .Q (n_1741));
  NA2X1 g63723(.A (n_6345), .B (csr_mcause_interrupt_flag), .Q
       (n_1739));
  NO2I1X1 g63724(.B (instruction[23]), .AN (instruction[22]), .Q
       (n_1738));
  NA2I1X2 g63725(.B (instruction[21]), .AN (n_1695), .Q (n_1737));
  NO2X1 g63726(.A (\instruction[8]_40015 ), .B (\instruction[7]_39562
       ), .Q (n_1736));
  NO2X1 g63727(.A (n_6603), .B (n_6600), .Q (n_1735));
  NO2I1X1 g63728(.B (csr_mcause_code[3]), .AN (csr_mcause_code[0]), .Q
       (n_1734));
  NO2X1 g63730(.A (csr_mcause_code[0]), .B (csr_mcause_code[3]), .Q
       (n_1733));
  NA2X1 g63731(.A (n_6453), .B (n_1688), .Q (n_1565));
  NO2I1X1 g63732(.B (csr_mcause_code[0]), .AN (csr_mcause_code[3]), .Q
       (n_1731));
  NA2I1X2 g63733(.B (n_1695), .AN (instruction[21]), .Q (n_1729));
  AND2X1 g63734(.A (csr_mcause_code[0]), .B (csr_mcause_code[3]), .Q
       (n_1728));
  NA2I1X4 g63735(.B (n_1578), .AN (instruction[23]), .Q (n_1582));
  NO2I1X1 g63736(.B (n_6720), .AN (n_6721), .Q (n_1727));
  NO2I1X1 g63737(.B (n_6721), .AN (n_6720), .Q (n_5606));
  NO2X1 g63738(.A (n_6601), .B (n_6604), .Q (jalr_type));
  NA2X4 g63739(.A (n_1580), .B (n_1694), .Q (n_1725));
  NA2X1 g63740(.A (n_6239), .B (n_1688), .Q (n_1723));
  NO2X1 g63741(.A (n_6071), .B (reset), .Q (n_1722));
  NO2X1 g63742(.A (n_1688), .B (reset), .Q (n_1721));
  NA2X4 g63743(.A (n_6720), .B (n_6721), .Q (n_1720));
  INX1 g63793(.A (n_6182), .Q (n_1714));
  INX1 g63794(.A (n_5146), .Q (n_1713));
  INX1 g63795(.A (n_5208), .Q (n_1712));
  INX1 g63796(.A (n_5351), .Q (n_1711));
  INX1 g63797(.A (n_5076), .Q (n_1710));
  INX1 g63798(.A (n_4979), .Q (n_1709));
  INX1 g63799(.A (n_4896), .Q (n_1708));
  INX1 g63800(.A (n_5204), .Q (n_1707));
  INX1 g63801(.A (n_4948), .Q (n_1706));
  INX1 g63802(.A (n_5201), .Q (n_1705));
  INX1 g63803(.A (n_4770), .Q (n_1704));
  INX1 g63804(.A (n_6010), .Q (n_1703));
  INX1 g63805(.A (n_6716), .Q (n_1702));
  INX1 g63807(.A (\instruction[11]_40800 ), .Q (n_1701));
  INX1 g63808(.A (\instruction[10]_39951 ), .Q (n_1700));
  INX1 g63809(.A (\instruction[9]_39983 ), .Q (n_1699));
  INX1 g63810(.A (system_type), .Q (n_1698));
  INX4 g63813(.A (flush_37507), .Q (n_6239));
  INX1 g63814(.A (n_4457), .Q (n_1697));
  INX1 g63815(.A (store_type), .Q (n_1696));
  BUX1 g63823(.A (n_6723), .Q (n_1695));
  INX4 g63824(.A (n_6723), .Q (n_1694));
  INX2 g63825(.A (n_6757), .Q (n_191));
  INX2 g63828(.A (instruction[24]), .Q (n_1690));
  INX1 g63829(.A (n_6459), .Q (n_1689));
  INX1 g63830(.A (n_6071), .Q (n_1688));
  INX1 g63832(.A (\instruction[5]_40139 ), .Q (n_1686));
  INX1 g63833(.A (n_5382), .Q (n_1685));
  INX1 g63834(.A (n_5212), .Q (n_1684));
  INX1 g63835(.A (n_5072), .Q (n_1683));
  INX1 g63836(.A (n_5320), .Q (n_1682));
  INX1 g63837(.A (n_4638), .Q (n_1681));
  INX1 g63838(.A (n_4895), .Q (n_1680));
  INX1 g63839(.A (n_5150), .Q (n_1679));
  INX1 g63840(.A (n_5134), .Q (n_1678));
  INX1 g63841(.A (n_4959), .Q (n_1677));
  INX1 g63842(.A (n_4961), .Q (n_1676));
  INX1 g63843(.A (n_5537), .Q (n_1675));
  INX1 g63844(.A (n_4607), .Q (n_1674));
  INX1 g63845(.A (n_4767), .Q (n_1673));
  INX1 g63846(.A (n_4762), .Q (n_1672));
  INX1 g63847(.A (n_5152), .Q (n_1671));
  INX1 g63848(.A (n_5103), .Q (n_1670));
  INX1 g63849(.A (n_5153), .Q (n_1669));
  INX1 g63850(.A (n_5475), .Q (n_1668));
  INX1 g63851(.A (n_5227), .Q (n_1667));
  INX1 g63852(.A (n_5413), .Q (n_1666));
  INX1 g63853(.A (n_5258), .Q (n_1665));
  INX1 g63854(.A (program_counter[2]), .Q (n_5574));
  INX1 g63855(.A (n_5542), .Q (n_1664));
  NA2I1X1 g41996(.B (n_1985), .AN (n_1574), .Q (n_1577));
  NA2I1X1 g63856(.B (n_1769), .AN (n_2997), .Q (n_1576));
  NA2I1X2 g63857(.B (n_1949), .AN (n_2081), .Q (n_1575));
  MU2IX2 g63858(.S (alu_operation_code_39061), .IN0 (n_177), .IN1
       (alu_2nd_operand[3]), .Q (n_6591));
  NA3I1X1 g63859(.B (n_1917), .C (n_3242), .AN (n_1975), .Q (n_1574));
  NA2I1X2 g63860(.B (n_1945), .AN (n_2077), .Q (n_1573));
  NO3I1X1 g63861(.B (n_1923), .C (n_3240), .AN (n_1912), .Q (n_1572));
  NA2I1X1 g63863(.B (n_2997), .AN (n_1769), .Q (n_1571));
  NA2I1X1 g63864(.B (n_1816), .AN (n_1770), .Q (n_1570));
  NA3I1X1 g63865(.B (csr_mcause_code[2]), .C (csr_mcause_code[4]), .AN
       (n_6373), .Q (n_1569));
  NO2I1X4 g63866(.B (n_1737), .AN (n_1839), .Q (n_1568));
  NO4I3X1 g63867(.D (csr_mcause_code[2]), .AN (n_1728), .BN (n_1802),
       .CN (csr_mcause_code[1]), .Q (irq_external_response));
  NA2I1X1 g63868(.B (n_1583), .AN (n_1582), .Q (n_1567));
  MU2X2 g63869(.S (n_1687), .IN0 (n_6014), .IN1 (\rs1_data[0]_39306 ),
       .Q (n_1566));
  NA2I1X1 g63872(.B (n_3037), .AN (n_4461), .Q (n_1564));
  INX1 g63876(.A (n_1594), .Q (n_1596));
  AND2X1 g63884(.A (n_2603), .B (n_2602), .Q (n_1616));
  AND2X1 g63886(.A (n_2745), .B (n_2738), .Q (n_1617));
  AND2X1 g63888(.A (n_2484), .B (n_2490), .Q (n_1611));
  AND2X1 g63890(.A (n_2470), .B (n_2464), .Q (n_1608));
  AND2X1 g63892(.A (n_2401), .B (n_2390), .Q (n_1605));
  AND2X1 g63894(.A (n_2414), .B (n_2402), .Q (n_1604));
  AND2X1 g63896(.A (n_2435), .B (n_2434), .Q (n_1609));
  AND2X1 g63898(.A (n_2431), .B (n_2432), .Q (n_1606));
  AND2X1 g63900(.A (n_2695), .B (n_2614), .Q (n_1614));
  AND2X1 g63902(.A (n_2703), .B (n_2621), .Q (n_1615));
  AND2X1 g63904(.A (n_2576), .B (n_2568), .Q (n_1619));
  AND2X1 g63906(.A (n_2555), .B (n_2556), .Q (n_1613));
  AND2X1 g63908(.A (n_2554), .B (n_2564), .Q (n_1612));
  AND2X1 g63910(.A (n_2739), .B (n_2751), .Q (n_1618));
  AND6X1 g63912(.A (n_2894), .B (n_2868), .C (n_2647), .D (n_2646), .E
       (n_2683), .F (n_2645), .Q (n_1630));
  AND6X1 g63914(.A (n_2889), .B (n_2873), .C (n_2665), .D (n_2664), .E
       (n_2690), .F (n_2663), .Q (n_1633));
  AND6X1 g63916(.A (n_2842), .B (n_2867), .C (n_2702), .D (n_2596), .E
       (n_2609), .F (n_2620), .Q (n_1626));
  AND6X1 g63918(.A (n_2828), .B (n_2825), .C (n_2567), .D (n_2531), .E
       (n_2494), .F (n_2495), .Q (n_1624));
  AND2X1 g63920(.A (n_2636), .B (n_2674), .Q (n_1620));
  INX1 g63924(.A (n_1589), .Q (n_1588));
  AND2X2 g63926(.A (n_1839), .B (n_1583), .Q (n_1590));
  INX2 g63928(.A (n_1947), .Q (n_1591));
  AND2X1 g63930(.A (instruction[21]), .B (n_1695), .Q (n_1583));
  AND2X1 g63932(.A (n_1727), .B (\instruction[14]_40077 ), .Q (n_6455));
  AND2X1 g63934(.A (n_6011), .B (n_1686), .Q (n_1581));
  OA21X1 g63936(.A (n_3100), .B (n_3093), .C (n_3099), .Q (n_1657));
  OA21X1 g63938(.A (n_6629), .B (n_6729), .C (n_3092), .Q (n_1654));
  OA21X1 g63940(.A (n_3122), .B (n_3096), .C (n_3121), .Q (n_1656));
  AND2X1 g63942(.A (n_1623), .B (n_1622), .Q (n_1643));
  AND2X1 g63944(.A (n_1634), .B (n_1629), .Q (n_1646));
  AND6X1 g63946(.A (n_1638), .B (n_2925), .C (n_2926), .D (n_2864), .E
       (n_2783), .F (n_2775), .Q (n_1648));
  AND6X1 g63948(.A (n_6746), .B (n_2817), .C (n_2529), .D (n_2527), .E
       (n_2528), .F (n_2519), .Q (n_1622));
  AND6X1 g63950(.A (n_2812), .B (n_2814), .C (n_2516), .D (n_2476), .E
       (n_2457), .F (n_2458), .Q (n_1621));
  AND6X1 g63952(.A (n_1614), .B (n_2840), .C (n_2696), .D (n_2708), .E
       (n_2697), .F (n_2615), .Q (n_1639));
  AND6X1 g63954(.A (n_2956), .B (n_2846), .C (n_2638), .D (n_2643), .E
       (n_2644), .F (n_2637), .Q (n_1627));
  AND6X1 g63956(.A (n_1615), .B (n_2853), .C (n_2704), .D (n_2709), .E
       (n_2622), .F (n_2613), .Q (n_1634));
  AND6X1 g63958(.A (n_2892), .B (n_2843), .C (n_2706), .D (n_2710), .E
       (n_2707), .F (n_2624), .Q (n_1640));
  AND6X1 g63960(.A (n_2887), .B (n_2871), .C (n_2659), .D (n_2658), .E
       (n_2688), .F (n_2657), .Q (n_1631));
  AND6X1 g63962(.A (n_6739), .B (n_2859), .C (n_2767), .D (n_2779), .E
       (n_2760), .F (n_2715), .Q (n_1636));
  AND6X1 g63964(.A (n_2951), .B (n_2865), .C (n_2774), .D (n_2729), .E
       (n_2676), .F (n_2678), .Q (n_1635));
  AND6X1 g63966(.A (n_1630), .B (n_2913), .C (n_2914), .D (n_2858), .E
       (n_2778), .F (n_2759), .Q (n_1650));
  AND6X1 g63968(.A (n_1633), .B (n_2928), .C (n_2906), .D (n_2955), .E
       (n_2785), .F (n_2764), .Q (n_1651));
  AND6X1 g63970(.A (n_1624), .B (n_2944), .C (n_2879), .D (n_2878), .E
       (n_2544), .F (n_2530), .Q (n_1645));
  AND6X1 g63972(.A (n_2835), .B (n_2826), .C (n_2551), .D (n_2552), .E
       (n_2553), .F (n_2563), .Q (n_1625));
  AND6X1 g63974(.A (n_2950), .B (n_2863), .C (n_2789), .D (n_2728), .E
       (n_2679), .F (n_2680), .Q (n_1642));
  AND6X1 g63976(.A (n_2948), .B (n_2945), .C (n_2790), .D (n_2755), .E
       (n_2712), .F (n_2711), .Q (n_1641));
  INX1 g63978(.A (n_211), .Q (n_5607));
  AND2X1 g63980(.A (n_1767), .B (n_1687), .Q (n_1586));
  AND2X1 g63982(.A (n_3105), .B (n_3108), .Q (n_1655));
  OA21X1 g63984(.A (n_3129), .B (n_3117), .C (n_3115), .Q (n_1658));
  AND6X1 g63986(.A (n_2821), .B (n_2811), .C (n_2487), .D (n_2485), .E
       (n_2492), .F (n_2486), .Q (n_1623));
  AND6X1 g63988(.A (n_1616), .B (n_6742), .C (n_2655), .D (n_2687), .E
       (n_2654), .F (n_2656), .Q (n_1629));
  AND6X1 g63990(.A (n_2910), .B (n_2949), .C (n_2743), .D (n_2747), .E
       (n_2742), .F (n_2753), .Q (n_1638));
  AND2X1 g63992(.A (n_1640), .B (n_1631), .Q (n_1647));
  AND6X1 g63994(.A (n_2893), .B (n_2869), .C (n_2649), .D (n_2684), .E
       (n_2685), .F (n_2648), .Q (n_1628));
  AND6X1 g63996(.A (n_1625), .B (n_2943), .C (n_2874), .D (n_2829), .E
       (n_2545), .F (n_2532), .Q (n_1644));
  AND6X1 g63998(.A (n_1642), .B (n_2942), .C (n_2924), .D (n_2934), .E
       (n_2746), .F (n_2741), .Q (n_1652));
  AND6X1 g64000(.A (n_1641), .B (n_2947), .C (n_2936), .D (n_2935), .E
       (n_2756), .F (n_2758), .Q (n_1653));
  OA21X1 g64002(.A (n_1662), .B (n_2084), .C (n_1799), .Q (n_1663));
  OA21X1 g64004(.A (n_3206), .B (n_3190), .C (n_3207), .Q (n_1660));
  AND6X1 g64006(.A (n_3191), .B (n_3189), .C (n_3193), .D (n_3171), .E
       (n_3169), .F (n_6725), .Q (n_1659));
  INX2 g64008(.A (n_1598), .Q (n_1599));
  AND6X1 g64010(.A (n_2927), .B (n_2866), .C (n_2776), .D (n_2784), .E
       (n_2763), .F (n_2732), .Q (n_1637));
  AND6X1 g64012(.A (n_2888), .B (n_2872), .C (n_2662), .D (n_2661), .E
       (n_2689), .F (n_2660), .Q (n_1632));
  OA21X1 g64014(.A (n_1714), .B (n_1934), .C (n_1986), .Q (n_204));
  OR3X2 g64016(.A (jalr_type), .B (store_type), .C (n_201), .Q
       (n_1587));
  AND6X1 g64018(.A (n_2983), .B (n_2979), .C (n_2911), .D (n_2890), .E
       (n_2899), .F (n_2898), .Q (n_1649));
  DFRQX1 \csr_mcause_reg[0] (.C (rc_gclk_205493), .D (n_693), .Q
       (csr_mcause[0]));
  DFRQX1 \csr_mcause_reg[10] (.C (rc_gclk_205493), .D (n_265), .Q
       (csr_mcause[10]));
  DFRQX1 \csr_mcause_reg[11] (.C (rc_gclk_205493), .D (n_104), .Q
       (csr_mcause[11]));
  DFRQX1 \csr_mcause_reg[12] (.C (rc_gclk_205493), .D (n_113), .Q
       (csr_mcause[12]));
  DFRQX1 \csr_mcause_reg[13] (.C (rc_gclk_205493), .D (n_103), .Q
       (csr_mcause[13]));
  DFRQX1 \csr_mcause_reg[14] (.C (rc_gclk_205493), .D (n_266), .Q
       (csr_mcause[14]));
  DFRQX1 \csr_mcause_reg[15] (.C (rc_gclk_205493), .D (n_102), .Q
       (csr_mcause[15]));
  DFRQX1 \csr_mcause_reg[16] (.C (rc_gclk_205493), .D (n_101), .Q
       (csr_mcause[16]));
  DFRQX1 \csr_mcause_reg[17] (.C (rc_gclk_205493), .D (n_100), .Q
       (csr_mcause[17]));
  DFRQX1 \csr_mcause_reg[18] (.C (rc_gclk_205493), .D (n_99), .Q
       (csr_mcause[18]));
  DFRQX1 \csr_mcause_reg[19] (.C (rc_gclk_205493), .D (n_98), .Q
       (csr_mcause[19]));
  DFRQX1 \csr_mcause_reg[1] (.C (rc_gclk_205493), .D (n_696), .Q
       (csr_mcause[1]));
  DFRQX1 \csr_mcause_reg[20] (.C (rc_gclk_205493), .D (n_258), .Q
       (csr_mcause[20]));
  DFRQX1 \csr_mcause_reg[21] (.C (rc_gclk_205493), .D (n_97), .Q
       (csr_mcause[21]));
  DFRQX1 \csr_mcause_reg[22] (.C (rc_gclk_205493), .D (n_112), .Q
       (csr_mcause[22]));
  DFRQX1 \csr_mcause_reg[23] (.C (rc_gclk_205493), .D (n_261), .Q
       (csr_mcause[23]));
  DFRQX1 \csr_mcause_reg[24] (.C (rc_gclk_205493), .D (n_96), .Q
       (csr_mcause[24]));
  DFRQX1 \csr_mcause_reg[25] (.C (rc_gclk_205493), .D (n_111), .Q
       (csr_mcause[25]));
  DFRQX1 \csr_mcause_reg[26] (.C (rc_gclk_205493), .D (n_110), .Q
       (csr_mcause[26]));
  DFRQX1 \csr_mcause_reg[27] (.C (rc_gclk_205493), .D (n_95), .Q
       (csr_mcause[27]));
  DFRQX1 \csr_mcause_reg[28] (.C (rc_gclk_205493), .D (n_109), .Q
       (csr_mcause[28]));
  DFRQX1 \csr_mcause_reg[29] (.C (rc_gclk_205493), .D (n_94), .Q
       (csr_mcause[29]));
  DFRQX1 \csr_mcause_reg[2] (.C (rc_gclk_205493), .D (n_710), .Q
       (csr_mcause[2]));
  DFRQX1 \csr_mcause_reg[30] (.C (rc_gclk_205493), .D (n_108), .Q
       (csr_mcause[30]));
  DFRQX1 \csr_mcause_reg[31] (.C (rc_gclk_205493), .D (n_694), .Q
       (csr_mcause[31]));
  DFRQX1 \csr_mcause_reg[3] (.C (rc_gclk_205493), .D (n_692), .Q
       (csr_mcause[3]));
  DFRQX1 \csr_mcause_reg[4] (.C (rc_gclk_205493), .D (n_695), .Q
       (csr_mcause[4]));
  DFRQX1 \csr_mcause_reg[5] (.C (rc_gclk_205493), .D (n_93), .Q
       (csr_mcause[5]));
  DFRQX1 \csr_mcause_reg[6] (.C (rc_gclk_205493), .D (n_92), .Q
       (csr_mcause[6]));
  DFRQX1 \csr_mcause_reg[7] (.C (rc_gclk_205493), .D (n_105), .Q
       (csr_mcause[7]));
  DFRQX1 \csr_mcause_reg[8] (.C (rc_gclk_205493), .D (n_107), .Q
       (csr_mcause[8]));
  DFRQX1 \csr_mcause_reg[9] (.C (rc_gclk_205493), .D (n_106), .Q
       (csr_mcause[9]));
  DFRQX1 \csr_mscratch_reg[0] (.C (rc_gclk_205577), .D (n_257), .Q
       (csr_mscratch[0]));
  DFRQX1 \csr_mscratch_reg[10] (.C (rc_gclk_205577), .D (n_91), .Q
       (csr_mscratch[10]));
  DFRQX1 \csr_mscratch_reg[11] (.C (rc_gclk_205577), .D (n_263), .Q
       (csr_mscratch[11]));
  DFRQX1 \csr_mscratch_reg[12] (.C (rc_gclk_205577), .D (n_113), .Q
       (csr_mscratch[12]));
  DFRQX1 \csr_mscratch_reg[13] (.C (rc_gclk_205577), .D (n_103), .Q
       (csr_mscratch[13]));
  DFRQX1 \csr_mscratch_reg[14] (.C (rc_gclk_205577), .D (n_90), .Q
       (csr_mscratch[14]));
  DFRQX1 \csr_mscratch_reg[15] (.C (rc_gclk_205577), .D (n_102), .Q
       (csr_mscratch[15]));
  DFRQX1 \csr_mscratch_reg[16] (.C (rc_gclk_205577), .D (n_101), .Q
       (csr_mscratch[16]));
  DFRQX1 \csr_mscratch_reg[17] (.C (rc_gclk_205577), .D (n_100), .Q
       (csr_mscratch[17]));
  DFRQX1 \csr_mscratch_reg[18] (.C (rc_gclk_205577), .D (n_264), .Q
       (csr_mscratch[18]));
  DFRQX1 \csr_mscratch_reg[19] (.C (rc_gclk_205577), .D (n_98), .Q
       (csr_mscratch[19]));
  DFRQX1 \csr_mscratch_reg[1] (.C (rc_gclk_205577), .D (n_406), .Q
       (csr_mscratch[1]));
  DFRQX1 \csr_mscratch_reg[20] (.C (rc_gclk_205577), .D (n_89), .Q
       (csr_mscratch[20]));
  DFRQX1 \csr_mscratch_reg[21] (.C (rc_gclk_205577), .D (n_259), .Q
       (csr_mscratch[21]));
  DFRQX1 \csr_mscratch_reg[22] (.C (rc_gclk_205577), .D (n_112), .Q
       (csr_mscratch[22]));
  DFRQX1 \csr_mscratch_reg[23] (.C (rc_gclk_205577), .D (n_88), .Q
       (csr_mscratch[23]));
  DFRQX1 \csr_mscratch_reg[24] (.C (rc_gclk_205577), .D (n_96), .Q
       (csr_mscratch[24]));
  DFRQX1 \csr_mscratch_reg[25] (.C (rc_gclk_205577), .D (n_111), .Q
       (csr_mscratch[25]));
  DFRQX1 \csr_mscratch_reg[26] (.C (rc_gclk_205577), .D (n_110), .Q
       (csr_mscratch[26]));
  DFRQX1 \csr_mscratch_reg[27] (.C (rc_gclk_205577), .D (n_262), .Q
       (csr_mscratch[27]));
  DFRQX1 \csr_mscratch_reg[28] (.C (rc_gclk_205577), .D (n_109), .Q
       (csr_mscratch[28]));
  DFRQX1 \csr_mscratch_reg[29] (.C (rc_gclk_205577), .D (n_267), .Q
       (csr_mscratch[29]));
  DFRQX1 \csr_mscratch_reg[2] (.C (rc_gclk_205577), .D (n_87), .Q
       (csr_mscratch[2]));
  DFRQX1 \csr_mscratch_reg[30] (.C (rc_gclk_205577), .D (n_108), .Q
       (csr_mscratch[30]));
  DFRQX1 \csr_mscratch_reg[31] (.C (rc_gclk_205577), .D (n_268), .Q
       (csr_mscratch[31]));
  DFRQX1 \csr_mscratch_reg[3] (.C (rc_gclk_205577), .D (n_86), .Q
       (csr_mscratch[3]));
  DFRQX1 \csr_mscratch_reg[4] (.C (rc_gclk_205577), .D (n_85), .Q
       (csr_mscratch[4]));
  DFRQX1 \csr_mscratch_reg[5] (.C (rc_gclk_205577), .D (n_254), .Q
       (csr_mscratch[5]));
  DFRQX1 \csr_mscratch_reg[6] (.C (rc_gclk_205577), .D (n_92), .Q
       (csr_mscratch[6]));
  DFRQX1 \csr_mscratch_reg[7] (.C (rc_gclk_205577), .D (n_105), .Q
       (csr_mscratch[7]));
  DFRQX1 \csr_mscratch_reg[8] (.C (rc_gclk_205577), .D (n_107), .Q
       (csr_mscratch[8]));
  DFRQX1 \csr_mscratch_reg[9] (.C (rc_gclk_205577), .D (n_106), .Q
       (csr_mscratch[9]));
  DFRQX1 csr_mstatus_mpie_reg(.C (rc_gclk), .D (n_939), .Q (n_4549));
  DFRQX1 \csr_mtval_reg[0] (.C (rc_gclk_205496), .D (n_868), .Q
       (csr_mtval[0]));
  DFRQX1 \csr_mtval_reg[10] (.C (rc_gclk_205496), .D (n_898), .Q
       (csr_mtval[10]));
  DFRQX1 \csr_mtval_reg[11] (.C (rc_gclk_205496), .D (n_902), .Q
       (csr_mtval[11]));
  DFRQX1 \csr_mtval_reg[12] (.C (rc_gclk_205496), .D (n_895), .Q
       (csr_mtval[12]));
  DFRQX1 \csr_mtval_reg[13] (.C (rc_gclk_205496), .D (n_894), .Q
       (csr_mtval[13]));
  DFRQX1 \csr_mtval_reg[14] (.C (rc_gclk_205496), .D (n_908), .Q
       (csr_mtval[14]));
  DFRQX1 \csr_mtval_reg[15] (.C (rc_gclk_205496), .D (n_907), .Q
       (csr_mtval[15]));
  DFRQX1 \csr_mtval_reg[16] (.C (rc_gclk_205496), .D (n_893), .Q
       (csr_mtval[16]));
  DFRQX1 \csr_mtval_reg[17] (.C (rc_gclk_205496), .D (n_892), .Q
       (csr_mtval[17]));
  DFRQX1 \csr_mtval_reg[18] (.C (rc_gclk_205496), .D (n_901), .Q
       (csr_mtval[18]));
  DFRQX1 \csr_mtval_reg[19] (.C (rc_gclk_205496), .D (n_897), .Q
       (csr_mtval[19]));
  DFRQX1 \csr_mtval_reg[1] (.C (rc_gclk_205496), .D (n_867), .Q
       (csr_mtval[1]));
  DFRQX1 \csr_mtval_reg[20] (.C (rc_gclk_205496), .D (n_896), .Q
       (csr_mtval[20]));
  DFRQX1 \csr_mtval_reg[21] (.C (rc_gclk_205496), .D (n_891), .Q
       (csr_mtval[21]));
  DFRQX1 \csr_mtval_reg[22] (.C (rc_gclk_205496), .D (n_903), .Q
       (csr_mtval[22]));
  DFRQX1 \csr_mtval_reg[23] (.C (rc_gclk_205496), .D (n_900), .Q
       (csr_mtval[23]));
  DFRQX1 \csr_mtval_reg[24] (.C (rc_gclk_205496), .D (n_890), .Q
       (csr_mtval[24]));
  DFRQX1 \csr_mtval_reg[25] (.C (rc_gclk_205496), .D (n_888), .Q
       (csr_mtval[25]));
  DFRQX1 \csr_mtval_reg[26] (.C (rc_gclk_205496), .D (n_906), .Q
       (csr_mtval[26]));
  DFRQX1 \csr_mtval_reg[27] (.C (rc_gclk_205496), .D (n_899), .Q
       (csr_mtval[27]));
  DFRQX1 \csr_mtval_reg[28] (.C (rc_gclk_205496), .D (n_909), .Q
       (csr_mtval[28]));
  DFRQX1 \csr_mtval_reg[29] (.C (rc_gclk_205496), .D (n_905), .Q
       (csr_mtval[29]));
  DFRQX1 \csr_mtval_reg[2] (.C (rc_gclk_205496), .D (n_886), .Q
       (csr_mtval[2]));
  DFRQX1 \csr_mtval_reg[30] (.C (rc_gclk_205496), .D (n_904), .Q
       (csr_mtval[30]));
  DFRQX1 \csr_mtval_reg[31] (.C (rc_gclk_205496), .D (n_911), .Q
       (csr_mtval[31]));
  DFRQX1 \csr_mtval_reg[3] (.C (rc_gclk_205496), .D (n_912), .Q
       (csr_mtval[3]));
  DFRQX1 \csr_mtval_reg[4] (.C (rc_gclk_205496), .D (n_910), .Q
       (csr_mtval[4]));
  DFRQX1 \csr_mtval_reg[5] (.C (rc_gclk_205496), .D (n_887), .Q
       (csr_mtval[5]));
  DFRQX1 \csr_mtval_reg[6] (.C (rc_gclk_205496), .D (n_889), .Q
       (csr_mtval[6]));
  DFRQX1 \csr_mtval_reg[7] (.C (rc_gclk_205496), .D (n_885), .Q
       (csr_mtval[7]));
  DFRQX1 \csr_mtval_reg[8] (.C (rc_gclk_205496), .D (n_862), .Q
       (csr_mtval[8]));
  DFRQX1 \csr_mtval_reg[9] (.C (rc_gclk_205496), .D (n_884), .Q
       (csr_mtval[9]));
  DFRQX1 \prev_instruction_address_reg[0] (.C (rc_gclk), .D (n_441), .Q
       (prev_instruction_address[0]));
  DFRQX1 \prev_instruction_address_reg[10] (.C (rc_gclk), .D (n_454),
       .Q (prev_instruction_address[10]));
  DFRQX1 \prev_instruction_address_reg[11] (.C (rc_gclk), .D (n_455),
       .Q (prev_instruction_address[11]));
  DFRQX1 \prev_instruction_address_reg[12] (.C (rc_gclk), .D (n_467),
       .Q (prev_instruction_address[12]));
  DFRQX1 \prev_instruction_address_reg[13] (.C (rc_gclk), .D (n_458),
       .Q (prev_instruction_address[13]));
  DFRQX1 \prev_instruction_address_reg[14] (.C (rc_gclk), .D (n_466),
       .Q (prev_instruction_address[14]));
  DFRQX1 \prev_instruction_address_reg[15] (.C (rc_gclk), .D (n_457),
       .Q (prev_instruction_address[15]));
  DFRQX1 \prev_instruction_address_reg[16] (.C (rc_gclk), .D (n_463),
       .Q (prev_instruction_address[16]));
  DFRQX1 \prev_instruction_address_reg[17] (.C (rc_gclk), .D (n_443),
       .Q (prev_instruction_address[17]));
  DFRQX1 \prev_instruction_address_reg[18] (.C (rc_gclk), .D (n_453),
       .Q (prev_instruction_address[18]));
  DFRQX1 \prev_instruction_address_reg[19] (.C (rc_gclk), .D (n_450),
       .Q (prev_instruction_address[19]));
  DFRQX1 \prev_instruction_address_reg[1] (.C (rc_gclk), .D (n_442), .Q
       (prev_instruction_address[1]));
  DFRQX1 \prev_instruction_address_reg[20] (.C (rc_gclk), .D (n_445),
       .Q (prev_instruction_address[20]));
  DFRQX1 \prev_instruction_address_reg[21] (.C (rc_gclk), .D (n_444),
       .Q (prev_instruction_address[21]));
  DFRQX1 \prev_instruction_address_reg[22] (.C (rc_gclk), .D (n_446),
       .Q (prev_instruction_address[22]));
  DFRQX1 \prev_instruction_address_reg[23] (.C (rc_gclk), .D (n_451),
       .Q (prev_instruction_address[23]));
  DFRQX1 \prev_instruction_address_reg[24] (.C (rc_gclk), .D (n_447),
       .Q (prev_instruction_address[24]));
  DFRQX1 \prev_instruction_address_reg[25] (.C (rc_gclk), .D (n_464),
       .Q (prev_instruction_address[25]));
  DFRQX1 \prev_instruction_address_reg[26] (.C (rc_gclk), .D (n_465),
       .Q (prev_instruction_address[26]));
  DFRQX1 \prev_instruction_address_reg[27] (.C (rc_gclk), .D (n_460),
       .Q (prev_instruction_address[27]));
  DFRQX1 \prev_instruction_address_reg[28] (.C (rc_gclk), .D (n_456),
       .Q (prev_instruction_address[28]));
  DFRQX1 \prev_instruction_address_reg[29] (.C (rc_gclk), .D (n_449),
       .Q (prev_instruction_address[29]));
  DFRQX1 \prev_instruction_address_reg[2] (.C (rc_gclk), .D (n_472), .Q
       (prev_instruction_address[2]));
  DFRQX1 \prev_instruction_address_reg[30] (.C (rc_gclk), .D (n_452),
       .Q (prev_instruction_address[30]));
  DFRQX1 \prev_instruction_address_reg[31] (.C (rc_gclk), .D (n_448),
       .Q (prev_instruction_address[31]));
  DFRQX1 \prev_instruction_address_reg[3] (.C (rc_gclk), .D (n_470), .Q
       (prev_instruction_address[3]));
  DFRQX1 \prev_instruction_address_reg[4] (.C (rc_gclk), .D (n_471), .Q
       (prev_instruction_address[4]));
  DFRQX1 \prev_instruction_address_reg[5] (.C (rc_gclk), .D (n_461), .Q
       (prev_instruction_address[5]));
  DFRQX1 \prev_instruction_address_reg[6] (.C (rc_gclk), .D (n_468), .Q
       (prev_instruction_address[6]));
  DFRQX1 \prev_instruction_address_reg[7] (.C (rc_gclk), .D (n_469), .Q
       (prev_instruction_address[7]));
  DFRQX1 \prev_instruction_address_reg[8] (.C (rc_gclk), .D (n_459), .Q
       (prev_instruction_address[8]));
  DFRQX1 \prev_instruction_address_reg[9] (.C (rc_gclk), .D (n_462), .Q
       (prev_instruction_address[9]));
  DFRQX1 \prev_instruction_reg[0] (.C (rc_gclk_205610), .D (n_239), .Q
       (prev_instruction[0]));
  DFRQX1 \prev_instruction_reg[10] (.C (rc_gclk_205610), .D (n_228), .Q
       (prev_instruction[10]));
  DFRQX1 \prev_instruction_reg[11] (.C (rc_gclk_205610), .D (n_227), .Q
       (prev_instruction[11]));
  DFRQX1 \prev_instruction_reg[12] (.C (rc_gclk_205610), .D (n_231), .Q
       (prev_instruction[12]));
  DFRQX1 \prev_instruction_reg[13] (.C (rc_gclk_205610), .D (n_233), .Q
       (prev_instruction[13]));
  DFRQX1 \prev_instruction_reg[14] (.C (rc_gclk_205610), .D (n_221), .Q
       (prev_instruction[14]));
  DFRQX1 \prev_instruction_reg[15] (.C (rc_gclk_205610), .D (n_251), .Q
       (prev_instruction[15]));
  DFRQX1 \prev_instruction_reg[16] (.C (rc_gclk_205610), .D (n_250), .Q
       (prev_instruction[16]));
  DFRQX1 \prev_instruction_reg[17] (.C (rc_gclk_205610), .D (n_252), .Q
       (prev_instruction[17]));
  DFRQX1 \prev_instruction_reg[18] (.C (rc_gclk_205610), .D (n_249), .Q
       (prev_instruction[18]));
  DFRQX1 \prev_instruction_reg[19] (.C (rc_gclk_205610), .D (n_246), .Q
       (prev_instruction[19]));
  DFRQX1 \prev_instruction_reg[1] (.C (rc_gclk_205610), .D (n_241), .Q
       (prev_instruction[1]));
  DFRQX1 \prev_instruction_reg[20] (.C (rc_gclk_205610), .D (n_248), .Q
       (prev_instruction[20]));
  DFRQX1 \prev_instruction_reg[21] (.C (rc_gclk_205610), .D (n_247), .Q
       (prev_instruction[21]));
  DFRQX1 \prev_instruction_reg[22] (.C (rc_gclk_205610), .D (n_244), .Q
       (prev_instruction[22]));
  DFRQX1 \prev_instruction_reg[23] (.C (rc_gclk_205610), .D (n_245), .Q
       (prev_instruction[23]));
  DFRQX1 \prev_instruction_reg[24] (.C (rc_gclk_205610), .D (n_243), .Q
       (prev_instruction[24]));
  DFRQX1 \prev_instruction_reg[25] (.C (rc_gclk_205610), .D (n_230), .Q
       (prev_instruction[25]));
  DFRQX1 \prev_instruction_reg[26] (.C (rc_gclk_205610), .D (n_225), .Q
       (prev_instruction[26]));
  DFRQX1 \prev_instruction_reg[27] (.C (rc_gclk_205610), .D (n_223), .Q
       (prev_instruction[27]));
  DFRQX1 \prev_instruction_reg[28] (.C (rc_gclk_205610), .D (n_220), .Q
       (prev_instruction[28]));
  DFRQX1 \prev_instruction_reg[29] (.C (rc_gclk_205610), .D (n_214), .Q
       (prev_instruction[29]));
  DFRQX1 \prev_instruction_reg[2] (.C (rc_gclk_205610), .D (n_238), .Q
       (prev_instruction[2]));
  DFRQX1 \prev_instruction_reg[30] (.C (rc_gclk_205610), .D (n_219), .Q
       (prev_instruction[30]));
  DFRQX1 \prev_instruction_reg[31] (.C (rc_gclk_205610), .D (n_218), .Q
       (prev_instruction[31]));
  DFRQX1 \prev_instruction_reg[3] (.C (rc_gclk_205610), .D (n_237), .Q
       (prev_instruction[3]));
  DFRQX1 \prev_instruction_reg[4] (.C (rc_gclk_205610), .D (n_240), .Q
       (prev_instruction[4]));
  DFRQX1 \prev_instruction_reg[5] (.C (rc_gclk_205610), .D (n_242), .Q
       (prev_instruction[5]));
  DFRQX1 \prev_instruction_reg[6] (.C (rc_gclk_205610), .D (n_234), .Q
       (prev_instruction[6]));
  DFRQX1 \prev_instruction_reg[7] (.C (rc_gclk_205610), .D (n_232), .Q
       (prev_instruction[7]));
  DFRQX1 \prev_instruction_reg[8] (.C (rc_gclk_205610), .D (n_216), .Q
       (prev_instruction[8]));
  DFRQX1 \prev_instruction_reg[9] (.C (rc_gclk_205610), .D (n_224), .Q
       (prev_instruction[9]));
  DFRQX1 \prev_rw_address_reg[0] (.C (rc_gclk), .D (n_477), .Q
       (prev_rw_address[0]));
  DFRQX1 \prev_rw_address_reg[10] (.C (rc_gclk), .D (n_499), .Q
       (prev_rw_address[10]));
  DFRQX1 \prev_rw_address_reg[11] (.C (rc_gclk), .D (n_502), .Q
       (prev_rw_address[11]));
  DFRQX1 \prev_rw_address_reg[12] (.C (rc_gclk), .D (n_506), .Q
       (prev_rw_address[12]));
  DFRQX1 \prev_rw_address_reg[13] (.C (rc_gclk), .D (n_504), .Q
       (prev_rw_address[13]));
  DFRQX1 \prev_rw_address_reg[14] (.C (rc_gclk), .D (n_503), .Q
       (prev_rw_address[14]));
  DFRQX1 \prev_rw_address_reg[15] (.C (rc_gclk), .D (n_501), .Q
       (prev_rw_address[15]));
  DFRQX1 \prev_rw_address_reg[16] (.C (rc_gclk), .D (n_507), .Q
       (prev_rw_address[16]));
  DFRQX1 \prev_rw_address_reg[17] (.C (rc_gclk), .D (n_486), .Q
       (prev_rw_address[17]));
  DFRQX1 \prev_rw_address_reg[18] (.C (rc_gclk), .D (n_493), .Q
       (prev_rw_address[18]));
  DFRQX1 \prev_rw_address_reg[19] (.C (rc_gclk), .D (n_485), .Q
       (prev_rw_address[19]));
  DFRQX1 \prev_rw_address_reg[1] (.C (rc_gclk), .D (n_495), .Q
       (prev_rw_address[1]));
  DFRQX1 \prev_rw_address_reg[20] (.C (rc_gclk), .D (n_487), .Q
       (prev_rw_address[20]));
  DFRQX1 \prev_rw_address_reg[21] (.C (rc_gclk), .D (n_494), .Q
       (prev_rw_address[21]));
  DFRQX1 \prev_rw_address_reg[22] (.C (rc_gclk), .D (n_492), .Q
       (prev_rw_address[22]));
  DFRQX1 \prev_rw_address_reg[23] (.C (rc_gclk), .D (n_489), .Q
       (prev_rw_address[23]));
  DFRQX1 \prev_rw_address_reg[24] (.C (rc_gclk), .D (n_488), .Q
       (prev_rw_address[24]));
  DFRQX1 \prev_rw_address_reg[25] (.C (rc_gclk), .D (n_505), .Q
       (prev_rw_address[25]));
  DFRQX1 \prev_rw_address_reg[26] (.C (rc_gclk), .D (n_498), .Q
       (prev_rw_address[26]));
  DFRQX1 \prev_rw_address_reg[27] (.C (rc_gclk), .D (n_490), .Q
       (prev_rw_address[27]));
  DFRQX1 \prev_rw_address_reg[28] (.C (rc_gclk), .D (n_508), .Q
       (prev_rw_address[28]));
  DFRQX1 \prev_rw_address_reg[29] (.C (rc_gclk), .D (n_491), .Q
       (prev_rw_address[29]));
  DFRQX1 \prev_rw_address_reg[2] (.C (rc_gclk), .D (n_481), .Q
       (prev_rw_address[2]));
  DFRQX1 \prev_rw_address_reg[30] (.C (rc_gclk), .D (n_483), .Q
       (prev_rw_address[30]));
  DFRQX1 \prev_rw_address_reg[31] (.C (rc_gclk), .D (n_484), .Q
       (prev_rw_address[31]));
  DFRQX1 \prev_rw_address_reg[3] (.C (rc_gclk), .D (n_479), .Q
       (prev_rw_address[3]));
  DFRQX1 \prev_rw_address_reg[4] (.C (rc_gclk), .D (n_482), .Q
       (prev_rw_address[4]));
  DFRQX1 \prev_rw_address_reg[5] (.C (rc_gclk), .D (n_500), .Q
       (prev_rw_address[5]));
  DFRQX1 \prev_rw_address_reg[6] (.C (rc_gclk), .D (n_480), .Q
       (prev_rw_address[6]));
  DFRQX1 \prev_rw_address_reg[7] (.C (rc_gclk), .D (n_478), .Q
       (prev_rw_address[7]));
  DFRQX1 \prev_rw_address_reg[8] (.C (rc_gclk), .D (n_496), .Q
       (prev_rw_address[8]));
  DFRQX1 \prev_rw_address_reg[9] (.C (rc_gclk), .D (n_497), .Q
       (prev_rw_address[9]));
  DFRQX1 \prev_write_data_reg[0] (.C (rc_gclk), .D (n_343), .Q
       (prev_write_data[0]));
  DFRQX1 \prev_write_data_reg[10] (.C (rc_gclk), .D (n_384), .Q
       (prev_write_data[10]));
  DFRQX1 \prev_write_data_reg[11] (.C (rc_gclk), .D (n_382), .Q
       (prev_write_data[11]));
  DFRQX1 \prev_write_data_reg[12] (.C (rc_gclk), .D (n_389), .Q
       (prev_write_data[12]));
  DFRQX1 \prev_write_data_reg[13] (.C (rc_gclk), .D (n_386), .Q
       (prev_write_data[13]));
  DFRQX1 \prev_write_data_reg[14] (.C (rc_gclk), .D (n_385), .Q
       (prev_write_data[14]));
  DFRQX1 \prev_write_data_reg[15] (.C (rc_gclk), .D (n_383), .Q
       (prev_write_data[15]));
  DFRQX1 \prev_write_data_reg[16] (.C (rc_gclk), .D (n_394), .Q
       (prev_write_data[16]));
  DFRQX1 \prev_write_data_reg[17] (.C (rc_gclk), .D (n_390), .Q
       (prev_write_data[17]));
  DFRQX1 \prev_write_data_reg[18] (.C (rc_gclk), .D (n_395), .Q
       (prev_write_data[18]));
  DFRQX1 \prev_write_data_reg[19] (.C (rc_gclk), .D (n_397), .Q
       (prev_write_data[19]));
  DFRQX1 \prev_write_data_reg[1] (.C (rc_gclk), .D (n_381), .Q
       (prev_write_data[1]));
  DFRQX1 \prev_write_data_reg[20] (.C (rc_gclk), .D (n_391), .Q
       (prev_write_data[20]));
  DFRQX1 \prev_write_data_reg[21] (.C (rc_gclk), .D (n_392), .Q
       (prev_write_data[21]));
  DFRQX1 \prev_write_data_reg[22] (.C (rc_gclk), .D (n_393), .Q
       (prev_write_data[22]));
  DFRQX1 \prev_write_data_reg[23] (.C (rc_gclk), .D (n_396), .Q
       (prev_write_data[23]));
  DFRQX1 \prev_write_data_reg[24] (.C (rc_gclk), .D (n_403), .Q
       (prev_write_data[24]));
  DFRQX1 \prev_write_data_reg[25] (.C (rc_gclk), .D (n_400), .Q
       (prev_write_data[25]));
  DFRQX1 \prev_write_data_reg[26] (.C (rc_gclk), .D (n_399), .Q
       (prev_write_data[26]));
  DFRQX1 \prev_write_data_reg[27] (.C (rc_gclk), .D (n_398), .Q
       (prev_write_data[27]));
  DFRQX1 \prev_write_data_reg[28] (.C (rc_gclk), .D (n_402), .Q
       (prev_write_data[28]));
  DFRQX1 \prev_write_data_reg[29] (.C (rc_gclk), .D (n_401), .Q
       (prev_write_data[29]));
  DFRQX1 \prev_write_data_reg[2] (.C (rc_gclk), .D (n_342), .Q
       (prev_write_data[2]));
  DFRQX1 \prev_write_data_reg[30] (.C (rc_gclk), .D (n_404), .Q
       (prev_write_data[30]));
  DFRQX1 \prev_write_data_reg[31] (.C (rc_gclk), .D (n_405), .Q
       (prev_write_data[31]));
  DFRQX1 \prev_write_data_reg[3] (.C (rc_gclk), .D (n_346), .Q
       (prev_write_data[3]));
  DFRQX1 \prev_write_data_reg[4] (.C (rc_gclk), .D (n_348), .Q
       (prev_write_data[4]));
  DFRQX1 \prev_write_data_reg[5] (.C (rc_gclk), .D (n_344), .Q
       (prev_write_data[5]));
  DFRQX1 \prev_write_data_reg[6] (.C (rc_gclk), .D (n_345), .Q
       (prev_write_data[6]));
  DFRQX1 \prev_write_data_reg[7] (.C (rc_gclk), .D (n_347), .Q
       (prev_write_data[7]));
  DFRQX1 \prev_write_data_reg[8] (.C (rc_gclk), .D (n_388), .Q
       (prev_write_data[8]));
  DFRQX1 \prev_write_data_reg[9] (.C (rc_gclk), .D (n_387), .Q
       (prev_write_data[9]));
  DFRQX1 \prev_write_strobe_reg[0] (.C (rc_gclk), .D (n_476), .Q
       (prev_write_strobe[0]));
  DFRQX1 \prev_write_strobe_reg[1] (.C (rc_gclk), .D (n_474), .Q
       (prev_write_strobe[1]));
  DFRQX1 \prev_write_strobe_reg[2] (.C (rc_gclk), .D (n_475), .Q
       (prev_write_strobe[2]));
  DFRQX1 \prev_write_strobe_reg[3] (.C (rc_gclk), .D (n_473), .Q
       (prev_write_strobe[3]));
  AN321X1 g47994(.A (n_119), .B (n_786), .C (n_1562), .D
       (program_counter[0]), .E (n_4532), .F (n_1527), .Q (n_1563));
  AN321X1 g47995(.A (n_878), .B (n_688), .C (n_1561), .D (n_858), .E
       (n_878), .F (n_1334), .Q (n_1562));
  AN32X1 g48680(.A (n_324), .B (n_339), .C (n_1548), .D (n_188), .E
       (alu_2nd_operand[15]), .Q (n_1561));
  AND3X1 g49346(.A (n_1054), .B (n_1481), .C (n_154), .Q (n_1560));
  AND3X1 g49347(.A (n_1068), .B (n_1418), .C (n_1536), .Q (n_1559));
  OA211X1 g49648(.A (n_1360), .B (n_970), .C (n_1448), .D (n_1544), .Q
       (n_1558));
  AND3X1 g49649(.A (n_1021), .B (n_1420), .C (n_1535), .Q (n_1557));
  ON22X1 g49877(.A (n_1528), .B (n_338), .C (n_210), .D
       (\rs1_data[14]_39466 ), .Q (n_1548));
  ON211X1 g49880(.A (n_1366), .B (n_977), .C (n_1524), .D (n_1423), .Q
       (n_1547));
  ON211X1 g49882(.A (n_1398), .B (n_968), .C (n_1388), .D (n_1521), .Q
       (n_1546));
  AND5X1 g49902(.A (n_1048), .B (n_1450), .C (n_567), .D (n_1461), .E
       (n_1489), .Q (n_1556));
  OA211X1 g49903(.A (n_1365), .B (n_970), .C (n_1447), .D (n_1520), .Q
       (n_1555));
  OA211X1 g49904(.A (n_1364), .B (n_970), .C (n_1537), .D (n_144), .Q
       (n_1554));
  OA211X1 g49905(.A (n_1367), .B (n_970), .C (n_1543), .D (n_141), .Q
       (n_1553));
  AND3X1 g49906(.A (n_1036), .B (n_1453), .C (n_1522), .Q (n_1552));
  AN21X1 g49907(.A (n_6078), .B (n_135), .C (n_1542), .Q (n_1551));
  OA211X1 g49908(.A (n_1371), .B (n_970), .C (n_1446), .D (n_1525), .Q
       (n_1550));
  AN21X1 g49909(.A (n_6073), .B (n_135), .C (n_1545), .Q (n_1549));
  ON211X1 g49939(.A (n_1359), .B (n_968), .C (n_1417), .D (n_1533), .Q
       (n_1545));
  AN21X1 g49951(.A (n_6085), .B (n_135), .C (n_1518), .Q (n_1544));
  AN21X1 g49953(.A (n_6082), .B (n_135), .C (n_1517), .Q (n_1543));
  ON211X1 g49954(.A (n_1361), .B (n_968), .C (n_1461), .D (n_1526), .Q
       (n_1542));
  ON211X1 g49955(.A (n_1371), .B (n_971), .C (n_1506), .D (n_1457), .Q
       (n_1541));
  ON211X1 g49956(.A (n_1357), .B (n_971), .C (n_1428), .D (n_1509), .Q
       (n_1540));
  ON211X1 g49957(.A (n_1367), .B (n_971), .C (n_1428), .D (n_1510), .Q
       (n_1539));
  NA3X1 g49958(.A (n_120), .B (n_1500), .C (n_1423), .Q (n_1538));
  AN21X1 g49960(.A (n_6083), .B (n_135), .C (n_1523), .Q (n_1537));
  AN211X1 g49961(.A (n_1002), .B (n_966), .C (n_1504), .D (n_1458), .Q
       (n_1536));
  AN221X1 g49962(.A (n_979), .B (n_991), .C (n_799), .D (read_data[6]),
       .E (n_1519), .Q (n_1535));
  ON211X1 g49963(.A (n_1213), .B (n_978), .C (n_142), .D (n_1502), .Q
       (n_1534));
  AN211X1 g49965(.A (n_5700), .B (n_270), .C (n_1488), .D (n_1458), .Q
       (n_1533));
  ON211X1 g49966(.A (n_1365), .B (n_971), .C (n_1429), .D (n_1497), .Q
       (n_1532));
  ON211X1 g49967(.A (n_1355), .B (n_977), .C (n_1423), .D (n_1498), .Q
       (n_1531));
  ON211X1 g49968(.A (n_1364), .B (n_971), .C (n_1429), .D (n_1516), .Q
       (n_1530));
  ON211X1 g49969(.A (n_1360), .B (n_971), .C (n_1457), .D (n_1496), .Q
       (n_1529));
  AN222X1 g49970(.A (n_193), .B (alu_2nd_operand[13]), .C (n_192), .D
       (alu_2nd_operand[12]), .E (n_1495), .F (n_938), .Q (n_1528));
  ON21X1 g49971(.A (n_1396), .B (n_970), .C (n_1505), .Q (n_1527));
  AN211X1 g49972(.A (n_5708), .B (n_270), .C (n_1494), .D (n_1297), .Q
       (n_1526));
  AND2X1 g49974(.A (n_1507), .B (n_1384), .Q (n_1525));
  AN21X1 g49975(.A (n_1004), .B (n_983), .C (n_1503), .Q (n_1524));
  NA3X1 g49976(.A (n_1348), .B (n_863), .C (n_1484), .Q (n_1523));
  AN211X1 g49977(.A (n_5709), .B (n_270), .C (n_1486), .D (n_1424), .Q
       (n_1522));
  AN221X1 g49978(.A (read_data[15]), .B (n_722), .C (n_1000), .D
       (n_966), .E (n_1490), .Q (n_1521));
  AN21X1 g49979(.A (n_799), .B (read_data[3]), .C (n_1501), .Q
       (n_1520));
  AO221X1 g49980(.A (n_270), .B (n_5711), .C (read_data[22]), .D
       (n_723), .E (n_1482), .Q (n_1519));
  AO211X1 g49981(.A (n_723), .B (read_data[18]), .C (n_796), .D
       (n_1485), .Q (n_1518));
  NA3X1 g49982(.A (n_1350), .B (n_950), .C (n_1483), .Q (n_1517));
  AN221X1 g49983(.A (n_985), .B (n_990), .C (n_1004), .D (n_979), .E
       (n_1472), .Q (n_1516));
  ON211X1 g49984(.A (n_1369), .B (n_977), .C (n_1478), .D (n_1456), .Q
       (n_1515));
  ON211X1 g49985(.A (n_1362), .B (n_977), .C (n_1423), .D (n_1479), .Q
       (n_1514));
  ON211X1 g49986(.A (n_1361), .B (n_977), .C (n_1480), .D (n_1455), .Q
       (n_1513));
  NA3X1 g49987(.A (n_1455), .B (n_1421), .C (n_1476), .Q (n_1512));
  ON211X1 g49988(.A (n_1449), .B (n_871), .C (n_1464), .D (n_882), .Q
       (n_1511));
  AN221X1 g49989(.A (n_985), .B (n_992), .C (n_996), .D (n_983), .E
       (n_1470), .Q (n_1510));
  AN221X1 g49990(.A (n_985), .B (n_991), .C (n_1013), .D (n_983), .E
       (n_1474), .Q (n_1509));
  NA3X1 g49991(.A (n_151), .B (n_1456), .C (n_1463), .Q (n_1508));
  AN221X1 g49992(.A (read_data[9]), .B (n_570), .C (n_723), .D
       (read_data[17]), .E (n_1465), .Q (n_1507));
  AN221X1 g49993(.A (n_961), .B (n_807), .C (n_997), .D (n_983), .E
       (n_1469), .Q (n_1506));
  AN211X1 g49994(.A (n_799), .B (read_data[0]), .C (n_1493), .D
       (n_1416), .Q (n_1505));
  ON221X1 g49996(.A (n_960), .B (n_806), .C (n_958), .D (n_814), .E
       (n_1499), .Q (n_1504));
  ON211X1 g49997(.A (n_846), .B (n_964), .C (n_1413), .D (n_1468), .Q
       (n_1503));
  AN221X1 g49998(.A (n_287), .B (n_729), .C (n_5710), .D (n_270), .E
       (n_1487), .Q (n_1502));
  ON211X1 g49999(.A (n_875), .B (n_962), .C (n_1466), .D (n_864), .Q
       (n_1501));
  AN221X1 g50000(.A (n_985), .B (n_1212), .C (n_1010), .D (n_979), .E
       (n_1475), .Q (n_1500));
  AN221X1 g50001(.A (read_data[13]), .B (n_722), .C (n_791), .D
       (n_1012), .E (n_1441), .Q (n_1499));
  NO3I1X1 g50002(.B (n_1345), .C (n_1343), .AN (n_1477), .Q (n_1498));
  AN21X1 g50003(.A (n_1011), .B (n_983), .C (n_1473), .Q (n_1497));
  AN21X1 g50004(.A (n_1003), .B (n_979), .C (n_1471), .Q (n_1496));
  ON311X1 g50005(.A (n_325), .B (n_326), .C (n_1452), .D (n_704), .E
       (n_663), .Q (n_1495));
  ON211X1 g50006(.A (n_806), .B (n_958), .C (n_1440), .D (n_1337), .Q
       (n_1494));
  NA2X1 g50007(.A (n_1335), .B (n_1467), .Q (n_1493));
  AN221X1 g50008(.A (read_data[12]), .B (n_722), .C (n_876), .D
       (n_1012), .E (n_1442), .Q (n_1492));
  ON221X1 g50009(.A (n_971), .B (n_1396), .C (n_871), .D (n_1351), .E
       (n_1445), .Q (n_1491));
  AO321X1 g50010(.A (n_874), .B (n_286), .C (n_581), .D
       (read_data[31]), .E (n_569), .F (n_1432), .Q (n_1490));
  AN221X1 g50011(.A (read_data[26]), .B (n_569), .C (n_722), .D
       (read_data[10]), .E (n_1433), .Q (n_1489));
  AO221X1 g50012(.A (read_data[14]), .B (n_722), .C (read_data[30]), .D
       (n_569), .E (n_1431), .Q (n_1488));
  AO221X1 g50013(.A (read_data[7]), .B (n_722), .C (read_data[23]), .D
       (n_569), .E (n_1434), .Q (n_1487));
  AO221X1 g50014(.A (read_data[8]), .B (n_722), .C (read_data[24]), .D
       (n_569), .E (n_1430), .Q (n_1486));
  ON211X1 g50015(.A (n_790), .B (n_962), .C (n_1437), .D (n_1444), .Q
       (n_1485));
  AN21X1 g50016(.A (n_5713), .B (n_270), .C (n_1462), .Q (n_1484));
  AN211X1 g50017(.A (n_571), .B (read_data[29]), .C (n_1438), .D
       (n_1427), .Q (n_1483));
  AO221X1 g50018(.A (read_data[14]), .B (n_570), .C (read_data[30]), .D
       (n_571), .E (n_1435), .Q (n_1482));
  AN21X1 g50019(.A (n_5705), .B (n_270), .C (n_1460), .Q (n_1481));
  AN211X1 g50020(.A (n_995), .B (n_980), .C (n_1410), .D (n_1390), .Q
       (n_1480));
  AN211X1 g50021(.A (n_989), .B (n_980), .C (n_1411), .D (n_1451), .Q
       (n_1479));
  AN221X1 g50022(.A (n_959), .B (n_791), .C (n_1349), .D (n_872), .E
       (n_1414), .Q (n_1478));
  AN221X1 g50023(.A (n_4483), .B (n_1148), .C (n_1214), .D (n_980), .E
       (n_1400), .Q (n_1477));
  AN221X1 g50024(.A (\rs1_data[26]_39276 ), .B (n_1152), .C (n_988), .D
       (n_980), .E (n_1406), .Q (n_1476));
  ON221X1 g50025(.A (n_981), .B (n_803), .C (n_982), .D (n_812), .E
       (n_145), .Q (n_1475));
  ON221X1 g50026(.A (n_962), .B (n_824), .C (n_964), .D (n_826), .E
       (n_146), .Q (n_1474));
  ON221X1 g50027(.A (n_962), .B (n_825), .C (n_964), .D (n_803), .E
       (n_149), .Q (n_1473));
  ON221X1 g50028(.A (n_981), .B (n_802), .C (n_982), .D (n_6764), .E
       (n_148), .Q (n_1472));
  ON221X1 g50029(.A (n_981), .B (n_828), .C (n_982), .D (n_821), .E
       (n_150), .Q (n_1471));
  ON221X1 g50030(.A (n_964), .B (n_808), .C (n_962), .D (n_822), .E
       (n_147), .Q (n_1470));
  ON21X1 g50031(.A (n_829), .B (n_964), .C (n_1436), .Q (n_1469));
  AN221X1 g50032(.A (\rs1_data[28]_39296 ), .B (n_1151), .C (n_876), .D
       (n_959), .E (n_1403), .Q (n_1468));
  AN221X1 g50033(.A (n_281), .B (n_994), .C (n_570), .D (read_data[8]),
       .E (n_1412), .Q (n_1467));
  AN211X1 g50034(.A (n_5714), .B (n_270), .C (n_1408), .D (n_1426), .Q
       (n_1466));
  NA2X1 g50035(.A (n_1444), .B (n_1439), .Q (n_1465));
  AN221X1 g50036(.A (n_133), .B (n_583), .C (n_987), .D (n_286), .E
       (n_1407), .Q (n_1464));
  AN221X1 g50037(.A (n_4485), .B (n_1150), .C (n_987), .D (n_576), .E
       (n_1401), .Q (n_1463));
  ON211X1 g50038(.A (n_319), .B (n_869), .C (n_1404), .D (n_1425), .Q
       (n_1462));
  INX1 g50039(.A (n_1459), .Q (n_1460));
  AN221X1 g50040(.A (n_984), .B (n_989), .C (n_1363), .D (n_967), .E
       (n_1393), .Q (n_1454));
  OA21X1 g50042(.A (n_1355), .B (n_968), .C (n_1419), .Q (n_1453));
  AN222X1 g50043(.A (n_187), .B (alu_2nd_operand[6]), .C (n_184), .D
       (alu_2nd_operand[5]), .E (n_1383), .F (n_327), .Q (n_1452));
  ON221X1 g50044(.A (n_981), .B (n_825), .C (n_982), .D (n_803), .E
       (n_1415), .Q (n_1451));
  AN221X1 g50045(.A (n_980), .B (n_1005), .C (n_1215), .D (n_967), .E
       (n_1391), .Q (n_1450));
  AN221X1 g50046(.A (n_282), .B (n_1010), .C (n_1397), .D
       (alu_2nd_operand[4]), .E (n_1336), .Q (n_1449));
  AN221X1 g50047(.A (read_data[2]), .B (n_799), .C (n_1005), .D
       (n_966), .E (n_1394), .Q (n_1448));
  AN221X1 g50048(.A (n_135), .B (n_6084), .C (n_998), .D (n_966), .E
       (n_1392), .Q (n_1447));
  AN211X1 g50049(.A (n_799), .B (read_data[1]), .C (n_1338), .D
       (n_1389), .Q (n_1446));
  AN211X1 g50050(.A (n_1324), .B (n_4484), .C (n_1377), .D (n_1395), .Q
       (n_1445));
  AN31X1 g50051(.A (alu_2nd_operand[4]), .B (alu_2nd_operand[1]), .C
       (n_1352), .D (n_1424), .Q (n_1461));
  AN21X1 g50052(.A (n_1352), .B (alu_2nd_operand[4]), .C (n_1424), .Q
       (n_1459));
  AO21X1 g50053(.A (n_1353), .B (n_294), .C (n_1424), .Q (n_1458));
  AN21X1 g50054(.A (n_1387), .B (alu_2nd_operand[1]), .C (n_1395), .Q
       (n_1457));
  NO2I1X1 g50055(.B (n_1353), .AN (n_1423), .Q (n_1456));
  AN21X1 g50056(.A (n_1352), .B (alu_2nd_operand[1]), .C (n_1422), .Q
       (n_1455));
  AN221X1 g50059(.A (n_4474), .B (n_1331), .C (n_569), .D
       (read_data[27]), .E (n_1379), .Q (n_1443));
  AO221X1 g50060(.A (read_data[28]), .B (n_569), .C
       (alu_2nd_operand[12]), .D (n_1308), .E (n_1373), .Q (n_1442));
  AO221X1 g50061(.A (read_data[29]), .B (n_569), .C
       (alu_2nd_operand[13]), .D (n_1307), .E (n_1372), .Q (n_1441));
  AN221X1 g50062(.A (n_4487), .B (n_1321), .C (n_569), .D
       (read_data[25]), .E (n_1375), .Q (n_1440));
  AN211X1 g50063(.A (n_5573), .B (n_270), .C (n_935), .D (n_1382), .Q
       (n_1439));
  ON21X1 g50064(.A (n_327), .B (n_869), .C (n_1399), .Q (n_1438));
  AN221X1 g50065(.A (n_6628), .B (n_1330), .C (n_5716), .D (n_270), .E
       (n_1378), .Q (n_1437));
  AN31X1 g50066(.A (n_872), .B (n_577), .C (n_581), .D (n_1409), .Q
       (n_1436));
  AO211X1 g50067(.A (n_1303), .B (alu_2nd_operand[6]), .C (n_1374), .D
       (n_1427), .Q (n_1435));
  AO211X1 g50068(.A (n_1302), .B (alu_2nd_operand[7]), .C (n_1385), .D
       (n_1386), .Q (n_1434));
  AO221X1 g50069(.A (n_4480), .B (n_1153), .C (n_1305), .D
       (alu_2nd_operand[10]), .E (n_6615), .Q (n_1433));
  ON211X1 g50070(.A (n_324), .B (n_869), .C (n_1354), .D (n_1402), .Q
       (n_1432));
  ON21X0 g50071(.A (n_339), .B (n_869), .C (n_1405), .Q (n_1431));
  AO221X1 g50072(.A (n_4464), .B (n_1147), .C (n_1298), .D
       (alu_2nd_operand[8]), .E (n_6614), .Q (n_1430));
  NA2X1 g50073(.A (n_1426), .B (alu_2nd_operand[1]), .Q (n_1444));
  INX1 g50074(.A (n_1425), .Q (n_1426));
  INX1 g50075(.A (n_1423), .Q (n_1422));
  AN221X1 g50076(.A (n_983), .B (n_1003), .C (n_1215), .D (n_976), .E
       (n_1339), .Q (n_1421));
  AN211X1 g50077(.A (n_1358), .B (n_969), .C (n_1344), .D (n_1346), .Q
       (n_1420));
  AN221X1 g50078(.A (n_984), .B (n_1214), .C (n_1009), .D (n_966), .E
       (n_1342), .Q (n_1419));
  AN22X1 g50079(.A (n_1370), .B (n_967), .C (n_5702), .D (n_270), .Q
       (n_1418));
  AN221X1 g50080(.A (n_957), .B (n_801), .C (n_999), .D (n_966), .E
       (n_1340), .Q (n_1417));
  ON221X1 g50081(.A (n_974), .B (n_816), .C (n_973), .D (n_809), .E
       (n_1376), .Q (n_1416));
  AN221X1 g50082(.A (n_961), .B (n_877), .C (n_834), .D (n_963), .E
       (n_1352), .Q (n_1415));
  ON221X1 g50083(.A (n_869), .B (n_545), .C (n_870), .D (n_235), .E
       (n_1326), .Q (n_1414));
  AN321X1 g50084(.A (n_4533), .B (\rs1_data[28]_39296 ), .C (n_994), .D
       (n_872), .E (n_856), .F (n_1352), .Q (n_1413));
  AO311X1 g50085(.A (n_866), .B (alu_sra_result[31]), .C (n_583), .D
       (n_928), .E (n_1332), .Q (n_1412));
  NO2X1 g50086(.A (n_1395), .B (n_1387), .Q (n_1429));
  AN21X1 g50087(.A (n_1353), .B (n_282), .C (n_1395), .Q (n_1428));
  NO2I1X1 g50088(.B (n_288), .AN (n_1386), .Q (n_1427));
  NA2X1 g50089(.A (n_1386), .B (alu_2nd_operand[2]), .Q (n_1425));
  OR2X1 g50090(.A (n_820), .B (n_1386), .Q (n_1424));
  NO2X1 g50091(.A (n_1395), .B (n_1368), .Q (n_1423));
  ON221X1 g50093(.A (n_194), .B (n_1329), .C (n_869), .D (n_304), .E
       (n_1320), .Q (n_1411));
  ON221X1 g50095(.A (n_199), .B (n_1323), .C (n_869), .D (n_311), .E
       (n_1314), .Q (n_1410));
  ON221X1 g50096(.A (n_869), .B (n_555), .C (n_870), .D (n_215), .E
       (n_1315), .Q (n_1409));
  AO221X1 g50098(.A (n_6757), .B (n_1325), .C (n_133), .D (n_328), .E
       (n_1317), .Q (n_1408));
  ON211X1 g50099(.A (n_236), .B (n_870), .C (n_1304), .D (n_1149), .Q
       (n_1407));
  AO221X1 g50101(.A (alu_2nd_operand[26]), .B (n_1312), .C (n_6453), .D
       (csr_data_out[26]), .E (n_926), .Q (n_1406));
  AN221X1 g50102(.A (n_134), .B (\rs1_data[14]_39466 ), .C (n_1313), .D
       (alu_2nd_operand[14]), .E (n_1142), .Q (n_1405));
  AN221X1 g50103(.A (n_134), .B (n_4465), .C (alu_2nd_operand[4]), .D
       (n_1301), .E (n_6617), .Q (n_1404));
  AO221X1 g50104(.A (alu_2nd_operand[28]), .B (n_1306), .C (n_6453), .D
       (csr_data_out[28]), .E (n_924), .Q (n_1403));
  AN221X1 g50105(.A (n_134), .B (\rs1_data[15]_39476 ), .C (n_1311), .D
       (alu_2nd_operand[15]), .E (n_1144), .Q (n_1402));
  AO221X1 g50106(.A (n_1300), .B (alu_2nd_operand[30]), .C (n_6453), .D
       (csr_data_out[30]), .E (n_921), .Q (n_1401));
  AO221X1 g50107(.A (alu_2nd_operand[24]), .B (n_1309), .C (n_6453), .D
       (csr_data_out[24]), .E (n_927), .Q (n_1400));
  AN221X1 g50108(.A (n_134), .B (n_4461), .C (n_1299), .D
       (alu_2nd_operand[5]), .E (n_6608), .Q (n_1399));
  INX1 g50109(.A (n_1397), .Q (n_1398));
  ON222X1 g50111(.A (n_648), .B (n_986), .C (n_958), .D (n_836), .E
       (n_993), .F (n_642), .Q (n_1394));
  ON221X1 g50112(.A (n_974), .B (n_805), .C (n_973), .D (n_6766), .E
       (n_1171), .Q (n_1393));
  ON222X1 g50114(.A (n_647), .B (n_986), .C (n_958), .D (n_842), .E
       (n_993), .F (n_643), .Q (n_1392));
  AO222X1 g50115(.A (n_975), .B (n_801), .C (n_984), .D (n_988), .E
       (n_972), .F (n_811), .Q (n_1391));
  ON221X1 g50116(.A (n_962), .B (n_830), .C (n_982), .D (n_829), .E
       (n_140), .Q (n_1390));
  ON321X1 g50120(.A (n_178), .B (n_293), .C (n_960), .D (n_974), .E
       (n_823), .F (n_1159), .Q (n_1389));
  AN221X1 g50121(.A (n_959), .B (n_819), .C (n_804), .D (n_957), .E
       (n_820), .Q (n_1388));
  ON222X1 g50122(.A (n_279), .B (n_803), .C (n_177), .D (n_1213), .E
       (n_812), .F (n_284), .Q (n_1397));
  MU2IX1 g50123(.S (alu_2nd_operand[3]), .IN0 (n_1009), .IN1 (n_1214),
       .Q (n_1396));
  NA2X1 g50124(.A (n_882), .B (n_1354), .Q (n_1395));
  AO221X1 g50125(.A (n_133), .B (n_325), .C (n_134), .D (n_4460), .E
       (n_6613), .Q (n_1385));
  AN222X1 g50126(.A (n_577), .B (n_994), .C (read_data[25]), .D
       (n_571), .E (n_6086), .F (n_135), .Q (n_1384));
  ON21X1 g50127(.A (n_180), .B (n_4465), .C (n_1333), .Q (n_1383));
  ON321X1 g50128(.A (n_136), .B (n_203), .C (n_179), .D (n_870), .E
       (n_256), .F (n_6611), .Q (n_1382));
  AND2X1 g50129(.A (n_1328), .B (n_925), .Q (n_1381));
  AND2X1 g50130(.A (n_1327), .B (n_923), .Q (n_1380));
  ON221X1 g50131(.A (n_869), .B (n_307), .C (n_870), .D (n_206), .E
       (n_6612), .Q (n_1379));
  ON221X0 g50132(.A (n_869), .B (n_115), .C (n_870), .D (n_124), .E
       (n_6609), .Q (n_1378));
  ON21X1 g50133(.A (n_340), .B (n_869), .C (n_1316), .Q (n_1377));
  OA222X1 g50134(.A (n_960), .B (n_687), .C (n_648), .D (n_993), .E
       (n_883), .F (n_958), .Q (n_1376));
  ON221X0 g50135(.A (n_869), .B (n_296), .C (n_870), .D (n_208), .E
       (n_6616), .Q (n_1375));
  AO221X1 g50136(.A (n_133), .B (n_326), .C (n_134), .D (n_4466), .E
       (n_6618), .Q (n_1374));
  ON221X1 g50137(.A (n_869), .B (n_337), .C (n_870), .D (n_192), .E
       (n_1143), .Q (n_1373));
  AO221X1 g50138(.A (n_133), .B (n_338), .C (n_134), .D (n_4476), .E
       (n_1141), .Q (n_1372));
  AND2X1 g50139(.A (n_1368), .B (alu_2nd_operand[2]), .Q (n_1387));
  NO2X1 g50140(.A (n_1354), .B (n_177), .Q (n_1386));
  INX1 g50141(.A (n_1369), .Q (n_1370));
  INX1 g50142(.A (n_1362), .Q (n_1363));
  INX1 g50143(.A (n_1357), .Q (n_1358));
  AN21X1 g50145(.A (n_1001), .B (n_282), .C (n_1209), .Q (n_1351));
  AN22X1 g50146(.A (n_992), .B (n_979), .C (n_799), .D (read_data[5]),
       .Q (n_1350));
  ON221X1 g50147(.A (n_580), .B (n_822), .C (n_579), .D (n_808), .E
       (n_1163), .Q (n_1349));
  AN22X1 g50148(.A (n_990), .B (n_979), .C (n_799), .D (read_data[4]),
       .Q (n_1348));
  AN221X1 g50149(.A (n_575), .B (n_880), .C (n_724), .D
       (\rs1_data[29]_39336 ), .E (n_865), .Q (n_1347));
  ON22X1 g50150(.A (n_818), .B (n_974), .C (n_800), .D (n_973), .Q
       (n_1346));
  ON22X1 g50152(.A (n_846), .B (n_962), .C (n_802), .D (n_982), .Q
       (n_1345));
  ON22X1 g50153(.A (n_836), .B (n_960), .C (n_840), .D (n_958), .Q
       (n_1344));
  ON22X1 g50154(.A (n_841), .B (n_964), .C (n_827), .D (n_981), .Q
       (n_1343));
  ON22X1 g50155(.A (n_816), .B (n_960), .C (n_809), .D (n_958), .Q
       (n_1342));
  AN22X1 g50158(.A (n_819), .B (n_975), .C (n_832), .D (n_957), .Q
       (n_1341));
  AO32X1 g50159(.A (n_874), .B (n_576), .C (n_581), .D (n_959), .E
       (n_817), .Q (n_1340));
  ON22X1 g50160(.A (n_824), .B (n_964), .C (n_881), .D (n_962), .Q
       (n_1339));
  ON22X1 g50161(.A (n_806), .B (n_973), .C (n_857), .D (n_873), .Q
       (n_1338));
  AN21X1 g50162(.A (n_722), .B (read_data[9]), .C (n_1162), .Q
       (n_1337));
  AO222X1 g50163(.A (n_573), .B (n_783), .C (n_575), .D (n_877), .E
       (n_4485), .F (n_724), .Q (n_1336));
  AN222X1 g50164(.A (n_135), .B (n_6087), .C (read_data[24]), .D
       (n_571), .E (n_723), .F (read_data[16]), .Q (n_1335));
  ON221X1 g50165(.A (n_859), .B (n_792), .C (n_730), .D (n_861), .E
       (n_860), .Q (n_1334));
  ON221X1 g50166(.A (n_328), .B (n_855), .C (n_191), .D
       (alu_2nd_operand[3]), .E (n_319), .Q (n_1333));
  ON211X1 g50167(.A (n_226), .B (n_870), .C (n_6619), .D (n_1154), .Q
       (n_1332));
  ON221X1 g50169(.A (n_136), .B (n_206), .C (n_869), .D
       (alu_2nd_operand[11]), .E (n_870), .Q (n_1331));
  ON221X1 g50170(.A (n_136), .B (n_124), .C (n_869), .D
       (alu_2nd_operand[2]), .E (n_870), .Q (n_1330));
  AN211X1 g50172(.A (alu_2nd_operand[27]), .B (n_137), .C (n_134), .D
       (n_919), .Q (n_1329));
  AN321X1 g50173(.A (n_4477), .B (n_137), .C (alu_2nd_operand[19]), .D
       (n_6453), .E (csr_data_out[19]), .F (n_920), .Q (n_1328));
  AN321X1 g50174(.A (n_4478), .B (n_137), .C (alu_2nd_operand[18]), .D
       (n_6453), .E (csr_data_out[18]), .F (n_913), .Q (n_1327));
  AN321X1 g50175(.A (\rs1_data[29]_39336 ), .B (n_137), .C
       (alu_2nd_operand[29]), .D (n_6453), .E (csr_data_out[29]), .F
       (n_922), .Q (n_1326));
  ON221X1 g50176(.A (n_136), .B (n_177), .C (n_869), .D
       (alu_2nd_operand[3]), .E (n_870), .Q (n_1325));
  ON211X1 g50177(.A (alu_2nd_operand[16]), .B (n_869), .C (n_870), .D
       (n_918), .Q (n_1324));
  AN211X1 g50178(.A (alu_2nd_operand[25]), .B (n_137), .C (n_134), .D
       (n_917), .Q (n_1323));
  AN321X1 g50179(.A (n_4486), .B (n_137), .C (alu_2nd_operand[20]), .D
       (n_6453), .E (csr_data_out[20]), .F (n_929), .Q (n_1322));
  ON221X1 g50180(.A (n_136), .B (n_208), .C (n_869), .D
       (alu_2nd_operand[9]), .E (n_870), .Q (n_1321));
  AN221X1 g50181(.A (n_6453), .B (csr_data_out[27]), .C
       (alu_2nd_operand[27]), .D (n_134), .E (n_934), .Q (n_1320));
  AN321X1 g50182(.A (n_4479), .B (n_137), .C (alu_2nd_operand[21]), .D
       (n_6453), .E (csr_data_out[21]), .F (n_930), .Q (n_1319));
  AN321X1 g50184(.A (n_4463), .B (n_137), .C (alu_2nd_operand[22]), .D
       (n_6453), .E (csr_data_out[22]), .F (n_931), .Q (n_1318));
  ON21X1 g50185(.A (n_177), .B (n_870), .C (n_6610), .Q (n_1317));
  AN221X1 g50186(.A (n_6453), .B (csr_data_out[16]), .C
       (alu_2nd_operand[16]), .D (n_134), .E (n_915), .Q (n_1316));
  AN321X1 g50187(.A (n_4482), .B (n_137), .C (alu_2nd_operand[17]), .D
       (n_6453), .E (csr_data_out[17]), .F (n_914), .Q (n_1315));
  AN221X1 g50188(.A (n_6453), .B (csr_data_out[25]), .C
       (alu_2nd_operand[25]), .D (n_134), .E (n_933), .Q (n_1314));
  ON221X1 g50189(.A (n_136), .B (n_197), .C (n_869), .D
       (\rs1_data[14]_39466 ), .E (n_870), .Q (n_1313));
  ON221X1 g50190(.A (n_136), .B (n_182), .C (n_869), .D
       (\rs1_data[26]_39276 ), .E (n_870), .Q (n_1312));
  ON221X1 g50191(.A (n_136), .B (n_188), .C (n_869), .D
       (\rs1_data[15]_39476 ), .E (n_870), .Q (n_1311));
  AN321X1 g50192(.A (\rs1_data[23]_39246 ), .B (n_137), .C
       (alu_2nd_operand[23]), .D (n_6453), .E (csr_data_out[23]), .F
       (n_932), .Q (n_1310));
  ON221X1 g50193(.A (n_136), .B (n_189), .C (n_869), .D (n_4483), .E
       (n_870), .Q (n_1309));
  ON221X1 g50194(.A (n_136), .B (n_192), .C (n_869), .D (n_4475), .E
       (n_870), .Q (n_1308));
  ON221X1 g50195(.A (n_136), .B (n_193), .C (n_869), .D (n_4476), .E
       (n_870), .Q (n_1307));
  ON221X1 g50196(.A (n_136), .B (n_181), .C (n_869), .D
       (\rs1_data[28]_39296 ), .E (n_870), .Q (n_1306));
  ON221X1 g50197(.A (n_136), .B (n_195), .C (n_869), .D (n_4480), .E
       (n_870), .Q (n_1305));
  AN211X1 g50198(.A (csr_data_out[31]), .B (n_6453), .C (n_936), .D
       (n_1210), .Q (n_1304));
  ON221X1 g50199(.A (n_136), .B (n_187), .C (n_869), .D (n_4466), .E
       (n_870), .Q (n_1303));
  ON221X1 g50200(.A (n_136), .B (n_196), .C (n_869), .D (n_4460), .E
       (n_870), .Q (n_1302));
  ON221X1 g50201(.A (n_136), .B (n_183), .C (n_869), .D (n_4465), .E
       (n_870), .Q (n_1301));
  ON221X1 g50202(.A (n_136), .B (n_186), .C (n_869), .D (n_4485), .E
       (n_870), .Q (n_1300));
  ON221X1 g50203(.A (n_136), .B (n_184), .C (n_869), .D (n_4461), .E
       (n_870), .Q (n_1299));
  ON221X1 g50204(.A (n_136), .B (n_190), .C (n_869), .D (n_4464), .E
       (n_870), .Q (n_1298));
  AO22X1 g50227(.A (n_1008), .B (n_966), .C (n_995), .D (n_984), .Q
       (n_1297));
  MU2IX1 g50228(.S (alu_2nd_operand[3]), .IN0 (n_1008), .IN1 (n_995),
       .Q (n_1371));
  MU2IX1 g50229(.S (alu_2nd_operand[3]), .IN0 (n_996), .IN1 (n_992), .Q
       (n_1369));
  NO2X1 g50230(.A (n_177), .B (n_1211), .Q (n_1368));
  AN22X1 g50231(.A (n_1002), .B (n_177), .C (n_791), .D (n_289), .Q
       (n_1367));
  AN21X1 g50232(.A (n_990), .B (alu_2nd_operand[3]), .C (n_952), .Q
       (n_1366));
  AN21X1 g50233(.A (n_989), .B (alu_2nd_operand[3]), .C (n_949), .Q
       (n_1365));
  AN22X1 g50234(.A (n_1007), .B (n_177), .C (n_876), .D (n_289), .Q
       (n_1364));
  AN21X1 g50235(.A (n_1011), .B (n_177), .C (n_943), .Q (n_1362));
  AN22X1 g50236(.A (n_997), .B (n_177), .C (n_582), .D (n_577), .Q
       (n_1361));
  AN222X1 g50237(.A (n_278), .B (n_801), .C (n_283), .D (n_811), .E
       (n_988), .F (alu_2nd_operand[3]), .Q (n_1360));
  MU2IX1 g50238(.S (alu_2nd_operand[3]), .IN0 (n_1013), .IN1 (n_991),
       .Q (n_1359));
  AN22X1 g50239(.A (n_999), .B (n_177), .C (n_582), .D (n_576), .Q
       (n_1357));
  AO22X1 g50240(.A (n_1000), .B (n_177), .C (n_582), .D (n_286), .Q
       (n_1356));
  AN22X1 g50241(.A (n_1001), .B (n_177), .C (n_582), .D (n_281), .Q
       (n_1355));
  NA2X1 g50242(.A (alu_2nd_operand[4]), .B (n_1210), .Q (n_1354));
  NO2X1 g50243(.A (n_288), .B (n_1211), .Q (n_1353));
  NO2X1 g50244(.A (n_284), .B (n_1211), .Q (n_1352));
  NO2X1 g50347(.A (n_1096), .B (n_123), .Q (n_1296));
  NO2X1 g50348(.A (n_1133), .B (n_123), .Q (n_1295));
  NO2X1 g50349(.A (n_1132), .B (n_123), .Q (n_1294));
  NO2X1 g50350(.A (n_1131), .B (n_123), .Q (n_1293));
  NO2X1 g50351(.A (n_1130), .B (n_123), .Q (n_1292));
  NO2X1 g50352(.A (n_1129), .B (n_123), .Q (n_1291));
  NO2X1 g50353(.A (n_1128), .B (n_123), .Q (n_1290));
  NO2X1 g50354(.A (n_1127), .B (n_123), .Q (n_1289));
  NO2X1 g50355(.A (n_1126), .B (n_123), .Q (n_1288));
  NO2X1 g50356(.A (n_1125), .B (n_123), .Q (n_1287));
  NO2X1 g50357(.A (n_1124), .B (n_123), .Q (n_1286));
  NO2X1 g50358(.A (n_1123), .B (n_123), .Q (n_1285));
  NO2X1 g50359(.A (n_1122), .B (n_123), .Q (n_1284));
  NO2X1 g50360(.A (n_1121), .B (n_123), .Q (n_1283));
  NO2X1 g50361(.A (n_1120), .B (n_123), .Q (n_1282));
  NO2X1 g50362(.A (n_1119), .B (n_123), .Q (n_1281));
  NO2X1 g50363(.A (n_1118), .B (n_123), .Q (n_1280));
  NO2X1 g50364(.A (n_1117), .B (n_123), .Q (n_1279));
  NO2X1 g50365(.A (n_1116), .B (n_123), .Q (n_1278));
  NO2X1 g50366(.A (n_1115), .B (n_123), .Q (n_1277));
  NO2X1 g50367(.A (n_1114), .B (n_123), .Q (n_1276));
  NO2X1 g50368(.A (n_1113), .B (n_123), .Q (n_1275));
  NO2X1 g50369(.A (n_1112), .B (n_123), .Q (n_1274));
  NO2X1 g50370(.A (n_1111), .B (n_123), .Q (n_1273));
  NO2X1 g50371(.A (n_1109), .B (n_123), .Q (n_1272));
  NO2X1 g50372(.A (n_1108), .B (n_123), .Q (n_1271));
  NO2X1 g50373(.A (n_1110), .B (n_123), .Q (n_1270));
  NO2X1 g50374(.A (n_1107), .B (n_123), .Q (n_1269));
  NO2X1 g50375(.A (n_1106), .B (n_123), .Q (n_1268));
  NO2X1 g50376(.A (n_1105), .B (n_123), .Q (n_1267));
  NO2X1 g50377(.A (n_1104), .B (n_123), .Q (n_1266));
  NO2X1 g50378(.A (n_1103), .B (n_123), .Q (n_1265));
  NO2X1 g50379(.A (n_1102), .B (n_123), .Q (n_1264));
  NO2X1 g50380(.A (n_1101), .B (n_123), .Q (n_1263));
  NO2X1 g50381(.A (n_1100), .B (n_123), .Q (n_1262));
  NO2X1 g50382(.A (n_1099), .B (n_123), .Q (n_1261));
  NO2X1 g50383(.A (n_1098), .B (n_123), .Q (n_1260));
  NO2X1 g50384(.A (n_1094), .B (n_123), .Q (n_1259));
  NO2X1 g50385(.A (n_1093), .B (n_123), .Q (n_1258));
  NO2X1 g50386(.A (n_1097), .B (n_123), .Q (n_1257));
  NO2X1 g50387(.A (n_1014), .B (n_123), .Q (n_1256));
  NO2X1 g50388(.A (n_1095), .B (n_123), .Q (n_1255));
  NO2X1 g50389(.A (n_1089), .B (n_123), .Q (n_1254));
  NO2X1 g50390(.A (n_1092), .B (n_123), .Q (n_1253));
  NO2X1 g50391(.A (n_1091), .B (n_123), .Q (n_1252));
  NO2X1 g50392(.A (n_1088), .B (n_123), .Q (n_1251));
  NO2X1 g50393(.A (n_1090), .B (n_123), .Q (n_1250));
  NO2X1 g50394(.A (n_1087), .B (n_123), .Q (n_1249));
  NO2X1 g50395(.A (n_1086), .B (n_123), .Q (n_1248));
  NO2X1 g50396(.A (n_1085), .B (n_123), .Q (n_1247));
  NO2X1 g50397(.A (n_1084), .B (n_123), .Q (n_1246));
  NO2X1 g50398(.A (n_1083), .B (n_123), .Q (n_1245));
  NO2X1 g50399(.A (n_1080), .B (n_123), .Q (n_1244));
  NO2X1 g50400(.A (n_1081), .B (n_123), .Q (n_1243));
  NO2X1 g50401(.A (n_1082), .B (n_123), .Q (n_1242));
  NO2X1 g50402(.A (n_1079), .B (n_123), .Q (n_1241));
  NO2X1 g50403(.A (n_1078), .B (n_123), .Q (n_1240));
  NO2X1 g50404(.A (n_1077), .B (n_123), .Q (n_1239));
  NO2X1 g50405(.A (n_1076), .B (n_123), .Q (n_1238));
  NO2X1 g50406(.A (n_1075), .B (n_123), .Q (n_1237));
  NO2X1 g50407(.A (n_1074), .B (n_123), .Q (n_1236));
  NO2X1 g50408(.A (n_1073), .B (n_123), .Q (n_1235));
  NO2X1 g50409(.A (n_1072), .B (n_123), .Q (n_1234));
  NO2X1 g50410(.A (n_1071), .B (n_123), .Q (n_1233));
  NO2X1 g50411(.A (n_1070), .B (n_123), .Q (n_1232));
  NO2X1 g50412(.A (n_1069), .B (n_123), .Q (n_1231));
  NO2X1 g50413(.A (n_1067), .B (n_123), .Q (n_1230));
  NO2X1 g50414(.A (n_1066), .B (n_123), .Q (n_1229));
  NO2X1 g50415(.A (n_1063), .B (n_123), .Q (n_1228));
  NO2X1 g50416(.A (n_1064), .B (n_123), .Q (n_1227));
  NO2X1 g50417(.A (n_1065), .B (n_123), .Q (n_1226));
  NO2X1 g50418(.A (n_1061), .B (n_123), .Q (n_1225));
  NO2X1 g50419(.A (n_1060), .B (n_123), .Q (n_1224));
  NO2X1 g50420(.A (n_1059), .B (n_123), .Q (n_1223));
  NO2X1 g50421(.A (n_1058), .B (n_123), .Q (n_1222));
  NO2X1 g50422(.A (n_1057), .B (n_123), .Q (n_1221));
  NO2X1 g50423(.A (n_1056), .B (n_123), .Q (n_1220));
  NO2X1 g50424(.A (n_1055), .B (n_123), .Q (n_1219));
  NO2X1 g50425(.A (n_1052), .B (n_123), .Q (n_1218));
  NO2X1 g50426(.A (n_1051), .B (n_123), .Q (n_1217));
  NO2X1 g50427(.A (n_1053), .B (n_123), .Q (n_1216));
  INX1 g50428(.A (n_1212), .Q (n_1213));
  INX1 g50429(.A (n_1211), .Q (n_1210));
  ON221X1 g50430(.A (n_574), .B (n_802), .C (n_572), .D (n_827), .E
       (n_691), .Q (n_1209));
  NO2X1 g50431(.A (n_1049), .B (n_123), .Q (n_1208));
  NO2X1 g50432(.A (n_1046), .B (n_123), .Q (n_1207));
  NO2X1 g50433(.A (n_1047), .B (n_123), .Q (n_1206));
  NO2X1 g50434(.A (n_1045), .B (n_123), .Q (n_1205));
  NO2X1 g50435(.A (n_1044), .B (n_123), .Q (n_1204));
  NO2X1 g50436(.A (n_1043), .B (n_123), .Q (n_1203));
  NO2X1 g50437(.A (n_1042), .B (n_123), .Q (n_1202));
  NO2X1 g50438(.A (n_1041), .B (n_123), .Q (n_1201));
  NO2X1 g50439(.A (n_1040), .B (n_123), .Q (n_1200));
  NO2X1 g50440(.A (n_1039), .B (n_123), .Q (n_1199));
  NO2X1 g50441(.A (n_1038), .B (n_123), .Q (n_1198));
  NO2X1 g50442(.A (n_1037), .B (n_123), .Q (n_1197));
  NO2X1 g50443(.A (n_1035), .B (n_123), .Q (n_1196));
  NO2X1 g50444(.A (n_1034), .B (n_123), .Q (n_1195));
  NO2X1 g50445(.A (n_1033), .B (n_123), .Q (n_1194));
  NO2X1 g50446(.A (n_1032), .B (n_123), .Q (n_1193));
  NO2X1 g50447(.A (n_1031), .B (n_123), .Q (n_1192));
  NO2X1 g50448(.A (n_1030), .B (n_123), .Q (n_1191));
  NO2X1 g50449(.A (n_1029), .B (n_123), .Q (n_1190));
  NO2X1 g50450(.A (n_1028), .B (n_123), .Q (n_1189));
  NO2X1 g50451(.A (n_1026), .B (n_123), .Q (n_1188));
  NO2X1 g50452(.A (n_1027), .B (n_123), .Q (n_1187));
  NO2X1 g50453(.A (n_1025), .B (n_123), .Q (n_1186));
  NO2X1 g50454(.A (n_1024), .B (n_123), .Q (n_1185));
  NO2X1 g50455(.A (n_1023), .B (n_123), .Q (n_1184));
  NO2X1 g50456(.A (n_1022), .B (n_123), .Q (n_1183));
  NO2X1 g50457(.A (n_1020), .B (n_123), .Q (n_1182));
  NO2X1 g50458(.A (n_1019), .B (n_123), .Q (n_1181));
  NO2X1 g50459(.A (n_1017), .B (n_123), .Q (n_1180));
  NO2X1 g50460(.A (n_1018), .B (n_123), .Q (n_1179));
  NO2X1 g50461(.A (n_1015), .B (n_123), .Q (n_1178));
  NO2X1 g50462(.A (n_1016), .B (n_123), .Q (n_1177));
  NO2X1 g50463(.A (n_1134), .B (n_123), .Q (n_1176));
  NO2X1 g50464(.A (n_951), .B (n_123), .Q (n_1175));
  NO2X1 g50465(.A (n_956), .B (n_123), .Q (n_1174));
  NO2X1 g50466(.A (n_955), .B (n_123), .Q (n_1173));
  NO2X1 g50467(.A (n_954), .B (n_123), .Q (n_1172));
  NA2X1 g50468(.A (n_998), .B (n_980), .Q (n_1171));
  NO2X1 g50469(.A (n_953), .B (n_123), .Q (n_1170));
  NO2X1 g50470(.A (n_1050), .B (n_123), .Q (n_1169));
  NO2X1 g50472(.A (n_948), .B (n_123), .Q (n_1167));
  NO2X1 g50473(.A (n_947), .B (n_123), .Q (n_1166));
  NO2X1 g50474(.A (n_946), .B (n_123), .Q (n_1165));
  AN221X1 g50476(.A (\rs1_data[28]_39296 ), .B (n_724), .C (n_831), .D
       (n_575), .E (n_853), .Q (n_1163));
  NO2X1 g50477(.A (n_823), .B (n_960), .Q (n_1162));
  NO2X1 g50478(.A (n_945), .B (n_123), .Q (n_1161));
  NO2X1 g50479(.A (n_944), .B (n_123), .Q (n_1160));
  OR2X1 g50480(.A (n_879), .B (n_958), .Q (n_1159));
  NO2X1 g50482(.A (n_942), .B (n_123), .Q (n_1157));
  NO2X1 g50483(.A (n_941), .B (n_123), .Q (n_1156));
  AND2X1 g50484(.A (n_937), .B (n_122), .Q (n_1155));
  AN22X1 g50485(.A (n_333), .B (n_137), .C (n_5604), .D (n_270), .Q
       (n_1154));
  ON21X1 g50486(.A (alu_2nd_operand[10]), .B (n_869), .C (n_870), .Q
       (n_1153));
  ON21X1 g50487(.A (alu_2nd_operand[26]), .B (n_869), .C (n_870), .Q
       (n_1152));
  ON21X1 g50488(.A (alu_2nd_operand[28]), .B (n_869), .C (n_870), .Q
       (n_1151));
  ON21X1 g50489(.A (alu_2nd_operand[30]), .B (n_869), .C (n_870), .Q
       (n_1150));
  NA3X1 g50490(.A (alu_2nd_operand[31]), .B (alu_sra_result[31]), .C
       (n_137), .Q (n_1149));
  ON21X1 g50491(.A (alu_2nd_operand[24]), .B (n_869), .C (n_870), .Q
       (n_1148));
  ON21X1 g50492(.A (alu_2nd_operand[8]), .B (n_869), .C (n_870), .Q
       (n_1147));
  AO222X1 g50495(.A (n_788), .B (n_6005), .C (n_6453), .D
       (csr_data_out[15]), .E (n_5587), .F (n_4532), .Q (n_1144));
  AN222X1 g50496(.A (n_788), .B (n_6008), .C (n_5584), .D (n_4532), .E
       (csr_data_out[12]), .F (n_6453), .Q (n_1143));
  AO222X1 g50497(.A (n_788), .B (n_6006), .C (n_6453), .D
       (csr_data_out[14]), .E (n_5586), .F (n_4532), .Q (n_1142));
  AO222X1 g50498(.A (n_788), .B (n_6007), .C (n_6453), .D
       (csr_data_out[13]), .E (n_5585), .F (n_4532), .Q (n_1141));
  ON222X1 g50505(.A (n_279), .B (n_828), .C (n_284), .D (n_821), .E
       (n_790), .F (n_290), .Q (n_1215));
  MU2X1 g50506(.S (alu_2nd_operand[2]), .IN0 (n_835), .IN1 (n_876), .Q
       (n_1214));
  MU2IX1 g50507(.S (n_124), .IN0 (n_875), .IN1 (n_793), .Q (n_1212));
  NA3X1 g50510(.A (alu_sra_result[31]), .B (n_874), .C
       (alu_operation_code_39061), .Q (n_1211));
  AN222X1 g50511(.A (n_5933), .B (n_131), .C (n_5934), .D (n_126), .E
       (n_5812), .F (n_125), .Q (n_1134));
  AN222X1 g50512(.A (n_131), .B (n_5819), .C (n_126), .D (n_5820), .E
       (n_5755), .F (n_125), .Q (n_1133));
  AN222X1 g50513(.A (n_131), .B (n_5827), .C (n_126), .D (n_5828), .E
       (n_5759), .F (n_125), .Q (n_1132));
  AN222X1 g50514(.A (n_117), .B (n_6303), .C (n_130), .D (n_6304), .E
       (n_6240), .F (n_129), .Q (n_1131));
  AN222X1 g50515(.A (n_117), .B (n_6305), .C (n_130), .D (n_6306), .E
       (n_6241), .F (n_129), .Q (n_1130));
  AN222X1 g50516(.A (n_117), .B (n_6311), .C (n_130), .D (n_6312), .E
       (n_6244), .F (n_129), .Q (n_1129));
  AN222X1 g50517(.A (n_131), .B (n_5823), .C (n_126), .D (n_5824), .E
       (n_5757), .F (n_125), .Q (n_1128));
  AN222X1 g50518(.A (n_117), .B (n_6307), .C (n_130), .D (n_6308), .E
       (n_6242), .F (n_129), .Q (n_1127));
  AN222X1 g50519(.A (n_131), .B (n_5829), .C (n_126), .D (n_5830), .E
       (n_5760), .F (n_125), .Q (n_1126));
  AN222X1 g50520(.A (n_131), .B (n_5835), .C (n_126), .D (n_5836), .E
       (n_5763), .F (n_125), .Q (n_1125));
  AN222X1 g50521(.A (n_117), .B (n_6313), .C (n_130), .D (n_6314), .E
       (n_6245), .F (n_129), .Q (n_1124));
  AN222X1 g50522(.A (n_117), .B (n_6319), .C (n_130), .D (n_6320), .E
       (n_6248), .F (n_129), .Q (n_1123));
  AN222X1 g50523(.A (n_131), .B (n_5825), .C (n_126), .D (n_5826), .E
       (n_5758), .F (n_125), .Q (n_1122));
  AN222X1 g50524(.A (n_131), .B (n_5831), .C (n_126), .D (n_5832), .E
       (n_5761), .F (n_125), .Q (n_1121));
  AN222X1 g50525(.A (n_131), .B (n_5851), .C (n_126), .D (n_5852), .E
       (n_5771), .F (n_125), .Q (n_1120));
  AN222X1 g50526(.A (n_131), .B (n_5843), .C (n_126), .D (n_5844), .E
       (n_5767), .F (n_125), .Q (n_1119));
  AN222X1 g50527(.A (n_131), .B (n_5837), .C (n_126), .D (n_5838), .E
       (n_5764), .F (n_125), .Q (n_1118));
  AN222X1 g50528(.A (n_117), .B (n_6309), .C (n_130), .D (n_6310), .E
       (n_6243), .F (n_129), .Q (n_1117));
  AN222X1 g50529(.A (n_117), .B (n_6315), .C (n_130), .D (n_6316), .E
       (n_6246), .F (n_129), .Q (n_1116));
  AN222X1 g50530(.A (n_131), .B (n_5833), .C (n_126), .D (n_5834), .E
       (n_5762), .F (n_125), .Q (n_1115));
  AN222X1 g50531(.A (n_117), .B (n_6357), .C (n_130), .D (n_6358), .E
       (n_6256), .F (n_129), .Q (n_1114));
  AN222X1 g50532(.A (n_117), .B (n_6349), .C (n_130), .D (n_6350), .E
       (n_6252), .F (n_129), .Q (n_1113));
  AN222X1 g50533(.A (n_117), .B (n_6321), .C (n_130), .D (n_6323), .E
       (n_6249), .F (n_129), .Q (n_1112));
  AN222X1 g50534(.A (n_117), .B (n_6317), .C (n_130), .D (n_6318), .E
       (n_6247), .F (n_129), .Q (n_1111));
  AN222X1 g50535(.A (n_131), .B (n_5845), .C (n_126), .D (n_5846), .E
       (n_5768), .F (n_125), .Q (n_1110));
  AN222X1 g50536(.A (n_131), .B (n_5859), .C (n_126), .D (n_5860), .E
       (n_5775), .F (n_125), .Q (n_1109));
  AN222X1 g50537(.A (n_131), .B (n_5853), .C (n_126), .D (n_5854), .E
       (n_5772), .F (n_125), .Q (n_1108));
  AN222X1 g50538(.A (n_131), .B (n_5839), .C (n_126), .D (n_5840), .E
       (n_5765), .F (n_125), .Q (n_1107));
  AN222X1 g50539(.A (n_117), .B (n_6365), .C (n_130), .D (n_6366), .E
       (n_6260), .F (n_129), .Q (n_1106));
  AN222X1 g50540(.A (n_117), .B (n_6359), .C (n_130), .D (n_6360), .E
       (n_6257), .F (n_129), .Q (n_1105));
  AN222X1 g50541(.A (n_117), .B (n_6351), .C (n_130), .D (n_6352), .E
       (n_6253), .F (n_129), .Q (n_1104));
  AN222X1 g50542(.A (n_117), .B (n_6329), .C (n_130), .D (n_6335), .E
       (n_6250), .F (n_129), .Q (n_1103));
  AN222X1 g50543(.A (n_131), .B (n_5867), .C (n_126), .D (n_5868), .E
       (n_5779), .F (n_125), .Q (n_1102));
  AN222X1 g50544(.A (n_131), .B (n_5861), .C (n_126), .D (n_5862), .E
       (n_5776), .F (n_125), .Q (n_1101));
  AN222X1 g50545(.A (n_131), .B (n_5855), .C (n_126), .D (n_5856), .E
       (n_5773), .F (n_125), .Q (n_1100));
  AN222X1 g50546(.A (n_131), .B (n_5847), .C (n_126), .D (n_5848), .E
       (n_5769), .F (n_125), .Q (n_1099));
  AN222X1 g50547(.A (n_131), .B (n_5841), .C (n_126), .D (n_5842), .E
       (n_5766), .F (n_125), .Q (n_1098));
  AN222X1 g50548(.A (n_117), .B (n_6375), .C (n_130), .D (n_6376), .E
       (n_6264), .F (n_129), .Q (n_1097));
  AN222X1 g50549(.A (n_117), .B (n_6368), .C (n_130), .D (n_6369), .E
       (n_6261), .F (n_129), .Q (n_1096));
  AN222X1 g50550(.A (n_117), .B (n_6361), .C (n_130), .D (n_6362), .E
       (n_6258), .F (n_129), .Q (n_1095));
  AN222X1 g50551(.A (n_117), .B (n_6353), .C (n_130), .D (n_6354), .E
       (n_6254), .F (n_129), .Q (n_1094));
  AN222X1 g50552(.A (n_117), .B (n_6341), .C (n_130), .D (n_6346), .E
       (n_6251), .F (n_129), .Q (n_1093));
  AN222X1 g50553(.A (n_131), .B (n_5857), .C (n_126), .D (n_5858), .E
       (n_5774), .F (n_125), .Q (n_1092));
  AN222X1 g50554(.A (n_131), .B (n_5875), .C (n_126), .D (n_5876), .E
       (n_5783), .F (n_125), .Q (n_1091));
  AN222X1 g50555(.A (n_131), .B (n_5869), .C (n_126), .D (n_5870), .E
       (n_5780), .F (n_125), .Q (n_1090));
  AN222X1 g50556(.A (n_131), .B (n_5863), .C (n_126), .D (n_5864), .E
       (n_5777), .F (n_125), .Q (n_1089));
  AN222X1 g50557(.A (n_131), .B (n_5849), .C (n_126), .D (n_5850), .E
       (n_5770), .F (n_125), .Q (n_1088));
  AN222X1 g50558(.A (n_117), .B (n_6383), .C (n_130), .D (n_6384), .E
       (n_6268), .F (n_129), .Q (n_1087));
  AN222X1 g50559(.A (n_117), .B (n_6377), .C (n_130), .D (n_6378), .E
       (n_6265), .F (n_129), .Q (n_1086));
  AN222X1 g50560(.A (n_117), .B (n_6370), .C (n_130), .D (n_6371), .E
       (n_6262), .F (n_129), .Q (n_1085));
  AN222X1 g50561(.A (n_117), .B (n_6363), .C (n_130), .D (n_6364), .E
       (n_6259), .F (n_129), .Q (n_1084));
  AN222X1 g50562(.A (n_117), .B (n_6355), .C (n_130), .D (n_6356), .E
       (n_6255), .F (n_129), .Q (n_1083));
  AN222X1 g50563(.A (n_131), .B (n_5877), .C (n_126), .D (n_5878), .E
       (n_5784), .F (n_125), .Q (n_1082));
  AN222X1 g50564(.A (n_131), .B (n_5871), .C (n_126), .D (n_5872), .E
       (n_5781), .F (n_125), .Q (n_1081));
  AN222X1 g50565(.A (n_131), .B (n_5865), .C (n_126), .D (n_5866), .E
       (n_5778), .F (n_125), .Q (n_1080));
  AN222X1 g50566(.A (n_117), .B (n_6385), .C (n_130), .D (n_6386), .E
       (n_6269), .F (n_129), .Q (n_1079));
  AN222X1 g50567(.A (n_117), .B (n_6379), .C (n_130), .D (n_6380), .E
       (n_6266), .F (n_129), .Q (n_1078));
  AN222X1 g50568(.A (n_117), .B (n_6372), .C (n_130), .D (n_6374), .E
       (n_6263), .F (n_129), .Q (n_1077));
  AN222X1 g50569(.A (n_131), .B (n_5879), .C (n_126), .D (n_5880), .E
       (n_5785), .F (n_125), .Q (n_1076));
  AN222X1 g50570(.A (n_131), .B (n_5873), .C (n_126), .D (n_5874), .E
       (n_5782), .F (n_125), .Q (n_1075));
  AN222X1 g50571(.A (n_6387), .B (n_117), .C (n_130), .D (n_6388), .E
       (n_6270), .F (n_129), .Q (n_1074));
  AN222X1 g50572(.A (n_6381), .B (n_117), .C (n_130), .D (n_6382), .E
       (n_6267), .F (n_129), .Q (n_1073));
  AN222X1 g50573(.A (n_131), .B (n_5881), .C (n_126), .D (n_5882), .E
       (n_5786), .F (n_125), .Q (n_1072));
  AN222X1 g50574(.A (n_6389), .B (n_117), .C (n_130), .D (n_6390), .E
       (n_6271), .F (n_129), .Q (n_1071));
  AN222X1 g50575(.A (n_131), .B (n_5883), .C (n_126), .D (n_5884), .E
       (n_5787), .F (n_125), .Q (n_1070));
  AN222X1 g50576(.A (n_6391), .B (n_117), .C (n_130), .D (n_6392), .E
       (n_6272), .F (n_129), .Q (n_1069));
  NA2X1 g50577(.A (n_6074), .B (n_135), .Q (n_1068));
  AN222X1 g50578(.A (n_131), .B (n_5885), .C (n_126), .D (n_5886), .E
       (n_5788), .F (n_125), .Q (n_1067));
  AN222X1 g50579(.A (n_131), .B (n_5891), .C (n_126), .D (n_5892), .E
       (n_5791), .F (n_125), .Q (n_1066));
  AN222X1 g50580(.A (n_6393), .B (n_117), .C (n_130), .D (n_6394), .E
       (n_6273), .F (n_129), .Q (n_1065));
  AN222X1 g50581(.A (n_6399), .B (n_117), .C (n_130), .D (n_6400), .E
       (n_6276), .F (n_129), .Q (n_1064));
  AN222X1 g50582(.A (n_6407), .B (n_117), .C (n_130), .D (n_6408), .E
       (n_6280), .F (n_129), .Q (n_1063));
  NA2X1 g50583(.A (n_6076), .B (n_135), .Q (n_1062));
  AN222X1 g50584(.A (n_131), .B (n_5887), .C (n_126), .D (n_5888), .E
       (n_5789), .F (n_125), .Q (n_1061));
  AN222X1 g50585(.A (n_131), .B (n_5907), .C (n_126), .D (n_5908), .E
       (n_5799), .F (n_125), .Q (n_1060));
  AN222X1 g50586(.A (n_131), .B (n_5893), .C (n_126), .D (n_5894), .E
       (n_5792), .F (n_125), .Q (n_1059));
  AN222X1 g50587(.A (n_6395), .B (n_117), .C (n_130), .D (n_6396), .E
       (n_6274), .F (n_129), .Q (n_1058));
  AN222X1 g50588(.A (n_6409), .B (n_117), .C (n_130), .D (n_6410), .E
       (n_6281), .F (n_129), .Q (n_1057));
  AN222X1 g50589(.A (n_6401), .B (n_117), .C (n_130), .D (n_6402), .E
       (n_6277), .F (n_129), .Q (n_1056));
  AN222X1 g50590(.A (n_6415), .B (n_117), .C (n_130), .D (n_6416), .E
       (n_6284), .F (n_129), .Q (n_1055));
  NA2X1 g50591(.A (n_6075), .B (n_135), .Q (n_1054));
  AN222X1 g50592(.A (n_5909), .B (n_131), .C (n_126), .D (n_5910), .E
       (n_5800), .F (n_125), .Q (n_1053));
  AN222X1 g50593(.A (n_5899), .B (n_131), .C (n_126), .D (n_5900), .E
       (n_5795), .F (n_125), .Q (n_1052));
  AN222X1 g50594(.A (n_5889), .B (n_131), .C (n_126), .D (n_5890), .E
       (n_5790), .F (n_125), .Q (n_1051));
  AN222X1 g50595(.A (n_5903), .B (n_131), .C (n_126), .D (n_5904), .E
       (n_5797), .F (n_125), .Q (n_1050));
  AN222X1 g50596(.A (n_5895), .B (n_131), .C (n_126), .D (n_5896), .E
       (n_5793), .F (n_125), .Q (n_1049));
  NA2X1 g50597(.A (n_6077), .B (n_135), .Q (n_1048));
  AN222X1 g50598(.A (n_6417), .B (n_117), .C (n_130), .D (n_6418), .E
       (n_6285), .F (n_129), .Q (n_1047));
  AN222X1 g50599(.A (n_6397), .B (n_117), .C (n_130), .D (n_6398), .E
       (n_6275), .F (n_129), .Q (n_1046));
  AN222X1 g50600(.A (n_6411), .B (n_117), .C (n_130), .D (n_6412), .E
       (n_6282), .F (n_129), .Q (n_1045));
  AN222X1 g50601(.A (n_6403), .B (n_117), .C (n_130), .D (n_6404), .E
       (n_6278), .F (n_129), .Q (n_1044));
  AN222X1 g50602(.A (n_5901), .B (n_131), .C (n_126), .D (n_5902), .E
       (n_5796), .F (n_125), .Q (n_1043));
  AN222X1 g50603(.A (n_5911), .B (n_131), .C (n_126), .D (n_5912), .E
       (n_5801), .F (n_125), .Q (n_1042));
  AN222X1 g50604(.A (n_5905), .B (n_131), .C (n_126), .D (n_5906), .E
       (n_5798), .F (n_125), .Q (n_1041));
  AN222X1 g50605(.A (n_5897), .B (n_131), .C (n_126), .D (n_5898), .E
       (n_5794), .F (n_125), .Q (n_1040));
  AN222X1 g50606(.A (n_6419), .B (n_117), .C (n_130), .D (n_6420), .E
       (n_6286), .F (n_129), .Q (n_1039));
  AN222X1 g50607(.A (n_6413), .B (n_117), .C (n_130), .D (n_6414), .E
       (n_6283), .F (n_129), .Q (n_1038));
  AN222X1 g50608(.A (n_6405), .B (n_117), .C (n_130), .D (n_6406), .E
       (n_6279), .F (n_129), .Q (n_1037));
  NA2X1 g50609(.A (n_6079), .B (n_135), .Q (n_1036));
  AN222X1 g50610(.A (n_5915), .B (n_131), .C (n_126), .D (n_5916), .E
       (n_5803), .F (n_125), .Q (n_1035));
  AN222X1 g50611(.A (n_5913), .B (n_131), .C (n_126), .D (n_5914), .E
       (n_5802), .F (n_125), .Q (n_1034));
  AN222X1 g50612(.A (n_6423), .B (n_117), .C (n_6424), .D (n_130), .E
       (n_6288), .F (n_129), .Q (n_1033));
  AN222X1 g50613(.A (n_6421), .B (n_117), .C (n_6422), .D (n_130), .E
       (n_6287), .F (n_129), .Q (n_1032));
  AN222X1 g50614(.A (n_5917), .B (n_131), .C (n_126), .D (n_5918), .E
       (n_5804), .F (n_125), .Q (n_1031));
  AN222X1 g50615(.A (n_5923), .B (n_131), .C (n_5924), .D (n_126), .E
       (n_5807), .F (n_125), .Q (n_1030));
  AN222X1 g50616(.A (n_6431), .B (n_117), .C (n_6432), .D (n_130), .E
       (n_6292), .F (n_129), .Q (n_1029));
  AN222X1 g50617(.A (n_6425), .B (n_117), .C (n_6426), .D (n_130), .E
       (n_6289), .F (n_129), .Q (n_1028));
  AN222X1 g50618(.A (n_5925), .B (n_131), .C (n_5926), .D (n_126), .E
       (n_5808), .F (n_125), .Q (n_1027));
  AN222X1 g50619(.A (n_5919), .B (n_131), .C (n_126), .D (n_5920), .E
       (n_5805), .F (n_125), .Q (n_1026));
  AN222X1 g50620(.A (n_6433), .B (n_117), .C (n_6434), .D (n_130), .E
       (n_6293), .F (n_129), .Q (n_1025));
  AN222X1 g50621(.A (n_6427), .B (n_117), .C (n_6428), .D (n_130), .E
       (n_6290), .F (n_129), .Q (n_1024));
  AN222X1 g50622(.A (n_5921), .B (n_131), .C (n_5922), .D (n_126), .E
       (n_5806), .F (n_125), .Q (n_1023));
  AN222X1 g50623(.A (n_5927), .B (n_131), .C (n_5928), .D (n_126), .E
       (n_5809), .F (n_125), .Q (n_1022));
  NA2X1 g50624(.A (n_6081), .B (n_135), .Q (n_1021));
  AN222X1 g50625(.A (n_6429), .B (n_117), .C (n_6430), .D (n_130), .E
       (n_6291), .F (n_129), .Q (n_1020));
  AN222X1 g50626(.A (n_6435), .B (n_117), .C (n_6436), .D (n_130), .E
       (n_6294), .F (n_129), .Q (n_1019));
  AN222X1 g50627(.A (n_5931), .B (n_131), .C (n_5932), .D (n_126), .E
       (n_5811), .F (n_125), .Q (n_1018));
  AN222X1 g50628(.A (n_5929), .B (n_131), .C (n_5930), .D (n_126), .E
       (n_5810), .F (n_125), .Q (n_1017));
  AN222X1 g50629(.A (n_6439), .B (n_117), .C (n_6440), .D (n_130), .E
       (n_6296), .F (n_129), .Q (n_1016));
  AN222X1 g50630(.A (n_6437), .B (n_117), .C (n_6438), .D (n_130), .E
       (n_6295), .F (n_129), .Q (n_1015));
  AN222X1 g50631(.A (n_131), .B (n_5821), .C (n_126), .D (n_5822), .E
       (n_5756), .F (n_125), .Q (n_1014));
  INX1 g50632(.A (n_1006), .Q (n_1007));
  INX1 g50633(.A (n_987), .Q (n_986));
  INX1 g50634(.A (n_979), .Q (n_978));
  INX1 g50635(.A (n_977), .Q (n_976));
  INX1 g50636(.A (n_975), .Q (n_974));
  INX1 g50637(.A (n_972), .Q (n_973));
  INX1 g50639(.A (n_970), .Q (n_969));
  INX1 g50640(.A (n_968), .Q (n_967));
  INX1 g50641(.A (n_966), .Q (n_965));
  INX1 g50642(.A (n_964), .Q (n_963));
  INX1 g50643(.A (n_962), .Q (n_961));
  INX1 g50644(.A (n_960), .Q (n_959));
  INX1 g50645(.A (n_958), .Q (n_957));
  AN222X1 g50647(.A (n_5935), .B (n_131), .C (n_5936), .D (n_126), .E
       (n_5813), .F (n_125), .Q (n_956));
  AN222X1 g50648(.A (n_6443), .B (n_117), .C (n_6444), .D (n_130), .E
       (n_6298), .F (n_129), .Q (n_955));
  AN222X1 g50649(.A (n_5937), .B (n_131), .C (n_5938), .D (n_126), .E
       (n_5814), .F (n_125), .Q (n_954));
  AN222X1 g50650(.A (n_5939), .B (n_131), .C (n_5940), .D (n_126), .E
       (n_5815), .F (n_125), .Q (n_953));
  ON22X1 g50651(.A (n_802), .B (n_279), .C (n_6764), .D (n_284), .Q
       (n_952));
  AN222X1 g50652(.A (n_6441), .B (n_117), .C (n_6442), .D (n_130), .E
       (n_6297), .F (n_129), .Q (n_951));
  AN222X0 g50654(.A (read_data[21]), .B (n_723), .C (read_data[13]), .D
       (n_570), .E (n_5712), .F (n_270), .Q (n_950));
  ON22X1 g50655(.A (n_805), .B (n_279), .C (n_6766), .D (n_284), .Q
       (n_949));
  AN222X1 g50666(.A (n_6445), .B (n_117), .C (n_6446), .D (n_130), .E
       (n_6299), .F (n_129), .Q (n_948));
  AN222X1 g50675(.A (n_6447), .B (n_117), .C (n_6448), .D (n_130), .E
       (n_6300), .F (n_129), .Q (n_947));
  AN222X1 g50678(.A (n_5941), .B (n_131), .C (n_5942), .D (n_126), .E
       (n_5816), .F (n_125), .Q (n_946));
  AN222X1 g50679(.A (n_6449), .B (n_117), .C (n_6450), .D (n_130), .E
       (n_6301), .F (n_129), .Q (n_945));
  AN222X1 g50680(.A (n_5943), .B (n_131), .C (n_5944), .D (n_126), .E
       (n_5817), .F (n_125), .Q (n_944));
  NO2X1 g50681(.A (n_875), .B (n_290), .Q (n_943));
  AN222X1 g50682(.A (n_5945), .B (n_131), .C (n_5946), .D (n_126), .E
       (n_5818), .F (n_125), .Q (n_942));
  AN222X1 g50683(.A (n_6451), .B (n_117), .C (n_6452), .D (n_130), .E
       (n_6302), .F (n_129), .Q (n_941));
  NO2X1 g50684(.A (n_854), .B (n_123), .Q (n_940));
  AO211X1 g50685(.A (n_6620), .B (n_4549), .C (n_123), .D (n_785), .Q
       (n_939));
  AN221X1 g50687(.A (n_705), .B (n_663), .C (n_554), .D (n_307), .E
       (n_336), .Q (n_938));
  ON22X1 g50690(.A (n_784), .B (csr_mcycle[0]), .C (n_4534), .D
       (n_568), .Q (n_937));
  AO222X1 g50698(.A (read_data[31]), .B (n_277), .C (n_6560), .D
       (n_788), .E (n_5603), .F (n_4532), .Q (n_936));
  AN21X1 g50699(.A (n_293), .B (n_334), .C (n_869), .Q (n_935));
  AO222X1 g50700(.A (read_data[27]), .B (n_277), .C (n_788), .D
       (n_5996), .E (n_5599), .F (n_4532), .Q (n_934));
  AO222X1 g50701(.A (read_data[25]), .B (n_277), .C (n_788), .D
       (n_5998), .E (n_5597), .F (n_4532), .Q (n_933));
  AO222X1 g50702(.A (read_data[23]), .B (n_277), .C (n_788), .D
       (n_6000), .E (n_5595), .F (n_4532), .Q (n_932));
  AO222X1 g50703(.A (read_data[22]), .B (n_277), .C (n_788), .D
       (n_5991), .E (n_5594), .F (n_4532), .Q (n_931));
  AO222X1 g50704(.A (read_data[21]), .B (n_277), .C (n_788), .D
       (n_6015), .E (n_5593), .F (n_4532), .Q (n_930));
  AO222X1 g50705(.A (read_data[20]), .B (n_277), .C (n_788), .D
       (n_5992), .E (n_5592), .F (n_4532), .Q (n_929));
  OA21X1 g50706(.A (n_281), .B (n_329), .C (n_133), .Q (n_928));
  AO222X1 g50707(.A (read_data[24]), .B (n_277), .C (n_788), .D
       (n_5999), .E (n_5596), .F (n_4532), .Q (n_927));
  AO222X1 g50708(.A (read_data[26]), .B (n_277), .C (n_788), .D
       (n_5997), .E (n_5598), .F (n_4532), .Q (n_926));
  ON21X1 g50709(.A (alu_2nd_operand[19]), .B (n_4477), .C (n_134), .Q
       (n_925));
  AO222X1 g50710(.A (read_data[28]), .B (n_277), .C (n_788), .D
       (n_5995), .E (n_5600), .F (n_4532), .Q (n_924));
  ON21X1 g50711(.A (alu_2nd_operand[18]), .B (n_4478), .C (n_134), .Q
       (n_923));
  AO222X1 g50712(.A (read_data[29]), .B (n_277), .C (n_788), .D
       (n_5994), .E (n_5601), .F (n_4532), .Q (n_922));
  AO222X1 g50713(.A (read_data[30]), .B (n_277), .C (n_788), .D
       (n_5993), .E (n_5602), .F (n_4532), .Q (n_921));
  AO222X1 g50714(.A (read_data[19]), .B (n_277), .C (n_788), .D
       (n_6001), .E (n_5591), .F (n_4532), .Q (n_920));
  NO2X1 g50715(.A (alu_2nd_operand[27]), .B (n_869), .Q (n_919));
  NA2X1 g50716(.A (alu_2nd_operand[16]), .B (n_137), .Q (n_918));
  NO2X1 g50717(.A (alu_2nd_operand[25]), .B (n_869), .Q (n_917));
  AO222X1 g50719(.A (read_data[16]), .B (n_277), .C (n_788), .D
       (n_6004), .E (n_5588), .F (n_4532), .Q (n_915));
  AO222X1 g50720(.A (read_data[17]), .B (n_277), .C (n_788), .D
       (n_6003), .E (n_5589), .F (n_4532), .Q (n_914));
  AO222X1 g50721(.A (read_data[18]), .B (n_277), .C (n_788), .D
       (n_6002), .E (n_5590), .F (n_4532), .Q (n_913));
  MU2IX1 g50722(.S (alu_2nd_operand[2]), .IN0 (n_845), .IN1 (n_828), .Q
       (n_1013));
  NO2X1 g50724(.A (n_655), .B (n_873), .Q (n_1012));
  MU2IX1 g50725(.S (alu_2nd_operand[2]), .IN0 (n_812), .IN1 (n_793), .Q
       (n_1011));
  MU2IX1 g50726(.S (alu_2nd_operand[2]), .IN0 (n_833), .IN1 (n_825), .Q
       (n_1010));
  MU2IX1 g50727(.S (alu_2nd_operand[2]), .IN0 (n_815), .IN1 (n_848), .Q
       (n_1009));
  MU2IX1 g50728(.S (alu_2nd_operand[2]), .IN0 (n_814), .IN1 (n_850), .Q
       (n_1008));
  MU2IX1 g50729(.S (alu_2nd_operand[2]), .IN0 (n_849), .IN1 (n_835), .Q
       (n_1006));
  MU2IX1 g50730(.S (alu_2nd_operand[2]), .IN0 (n_840), .IN1 (n_818), .Q
       (n_1005));
  MU2IX1 g50731(.S (alu_2nd_operand[2]), .IN0 (n_841), .IN1 (n_827), .Q
       (n_1004));
  MU2IX1 g50732(.S (alu_2nd_operand[2]), .IN0 (n_826), .IN1 (n_845), .Q
       (n_1003));
  MU2IX1 g50733(.S (alu_2nd_operand[2]), .IN0 (n_850), .IN1 (n_844), .Q
       (n_1002));
  MU2IX1 g50734(.S (alu_2nd_operand[2]), .IN0 (n_6764), .IN1 (n_132),
       .Q (n_1001));
  MU2IX1 g50735(.S (alu_2nd_operand[2]), .IN0 (n_6766), .IN1 (n_839),
       .Q (n_1000));
  MU2X1 g50736(.S (n_124), .IN0 (n_837), .IN1 (n_811), .Q (n_999));
  MU2X1 g50737(.S (alu_2nd_operand[2]), .IN0 (n_832), .IN1 (n_819), .Q
       (n_998));
  MU2IX1 g50738(.S (alu_2nd_operand[2]), .IN0 (n_6762), .IN1 (n_852),
       .Q (n_997));
  MU2IX1 g50739(.S (alu_2nd_operand[2]), .IN0 (n_829), .IN1 (n_6762),
       .Q (n_996));
  MU2X1 g50740(.S (alu_2nd_operand[2]), .IN0 (n_843), .IN1 (n_791), .Q
       (n_995));
  NO2X1 g50741(.A (n_578), .B (n_871), .Q (n_994));
  NA2X1 g50742(.A (n_726), .B (n_874), .Q (n_993));
  AO22X1 g50743(.A (n_851), .B (n_124), .C (n_292), .D (n_577), .Q
       (n_992));
  MU2IX1 g50744(.S (alu_2nd_operand[2]), .IN0 (n_821), .IN1 (n_790), .Q
       (n_991));
  ON22X1 g50745(.A (n_132), .B (alu_2nd_operand[2]), .C (n_291), .D
       (n_280), .Q (n_990));
  AO22X1 g50746(.A (n_838), .B (n_124), .C (n_292), .D (n_286), .Q
       (n_989));
  AO22X1 g50747(.A (n_837), .B (n_124), .C (n_292), .D (n_576), .Q
       (n_988));
  NO2X1 g50748(.A (n_578), .B (n_873), .Q (n_987));
  AND2X1 g50749(.A (n_294), .B (n_872), .Q (n_985));
  AND2X1 g50750(.A (n_294), .B (n_874), .Q (n_984));
  AND2X1 g50751(.A (n_282), .B (n_872), .Q (n_983));
  OR2X1 g50752(.A (n_579), .B (n_871), .Q (n_982));
  OR2X1 g50753(.A (n_580), .B (n_871), .Q (n_981));
  AND2X1 g50754(.A (n_310), .B (n_874), .Q (n_980));
  AND2X1 g50755(.A (n_310), .B (n_872), .Q (n_979));
  NA2X1 g50756(.A (alu_2nd_operand[4]), .B (n_872), .Q (n_977));
  NO2X1 g50757(.A (n_580), .B (n_873), .Q (n_975));
  NO2X1 g50758(.A (n_579), .B (n_873), .Q (n_972));
  NA2X1 g50759(.A (n_180), .B (n_874), .Q (n_971));
  NA2X1 g50760(.A (alu_2nd_operand[4]), .B (n_874), .Q (n_970));
  NA2X1 g50761(.A (n_180), .B (n_872), .Q (n_968));
  AND2X1 g50762(.A (n_282), .B (n_874), .Q (n_966));
  NA2X1 g50763(.A (n_575), .B (n_872), .Q (n_964));
  NA2X1 g50764(.A (n_573), .B (n_872), .Q (n_962));
  NA2X1 g50765(.A (n_573), .B (n_874), .Q (n_960));
  NA2X1 g50766(.A (n_575), .B (n_874), .Q (n_958));
  AN21X1 g50767(.A (n_532), .B (n_714), .C (n_123), .Q (n_912));
  AN21X1 g50768(.A (n_510), .B (n_715), .C (n_123), .Q (n_911));
  AN21X1 g50769(.A (n_533), .B (n_712), .C (n_123), .Q (n_910));
  AN21X1 g50770(.A (n_528), .B (n_720), .C (n_123), .Q (n_909));
  AN21X1 g50771(.A (n_514), .B (n_738), .C (n_123), .Q (n_908));
  AN21X1 g50772(.A (n_515), .B (n_748), .C (n_123), .Q (n_907));
  AN21X1 g50773(.A (n_526), .B (n_746), .C (n_123), .Q (n_906));
  AN21X1 g50774(.A (n_529), .B (n_718), .C (n_123), .Q (n_905));
  AN21X1 g50775(.A (n_531), .B (n_716), .C (n_123), .Q (n_904));
  AN21X1 g50776(.A (n_522), .B (n_732), .C (n_123), .Q (n_903));
  AN21X1 g50777(.A (n_511), .B (n_740), .C (n_123), .Q (n_902));
  AN21X1 g50778(.A (n_518), .B (n_736), .C (n_123), .Q (n_901));
  AN21X1 g50779(.A (n_523), .B (n_731), .C (n_123), .Q (n_900));
  AN21X1 g50780(.A (n_527), .B (n_719), .C (n_123), .Q (n_899));
  AN21X1 g50781(.A (n_539), .B (n_711), .C (n_123), .Q (n_898));
  AN21X1 g50782(.A (n_519), .B (n_735), .C (n_123), .Q (n_897));
  AN21X1 g50783(.A (n_520), .B (n_745), .C (n_123), .Q (n_896));
  AN21X1 g50784(.A (n_512), .B (n_749), .C (n_123), .Q (n_895));
  AN21X1 g50785(.A (n_513), .B (n_739), .C (n_123), .Q (n_894));
  AN21X1 g50786(.A (n_516), .B (n_737), .C (n_123), .Q (n_893));
  AN21X1 g50787(.A (n_517), .B (n_747), .C (n_123), .Q (n_892));
  AN21X1 g50788(.A (n_521), .B (n_733), .C (n_123), .Q (n_891));
  AN21X1 g50789(.A (n_524), .B (n_721), .C (n_123), .Q (n_890));
  AN21X1 g50790(.A (n_535), .B (n_742), .C (n_123), .Q (n_889));
  AN21X1 g50791(.A (n_525), .B (n_744), .C (n_123), .Q (n_888));
  AN21X1 g50792(.A (n_534), .B (n_734), .C (n_123), .Q (n_887));
  AN21X1 g50793(.A (n_530), .B (n_717), .C (n_123), .Q (n_886));
  AN21X1 g50794(.A (n_536), .B (n_741), .C (n_123), .Q (n_885));
  AN21X1 g50795(.A (n_537), .B (n_713), .C (n_123), .Q (n_884));
  INX1 g50796(.A (n_880), .Q (n_881));
  INX1 g50797(.A (n_874), .Q (n_873));
  INX1 g50798(.A (n_872), .Q (n_871));
  NO2X1 g50802(.A (n_795), .B (n_123), .Q (n_868));
  NO2X1 g50803(.A (n_794), .B (n_123), .Q (n_867));
  NO2X1 g50804(.A (n_789), .B (n_6597), .Q (n_866));
  NO2X1 g50805(.A (n_824), .B (n_580), .Q (n_865));
  AN222X1 g50806(.A (read_data[27]), .B (n_571), .C (read_data[11]), .D
       (n_570), .E (n_723), .F (read_data[19]), .Q (n_864));
  AN222X1 g50807(.A (read_data[28]), .B (n_571), .C (read_data[12]), .D
       (n_570), .E (n_723), .F (read_data[20]), .Q (n_863));
  AN21X1 g50808(.A (n_538), .B (n_743), .C (n_123), .Q (n_862));
  AN22X1 g50809(.A (n_661), .B (n_689), .C (n_553), .D (n_304), .Q
       (n_861));
  AN22X1 g50810(.A (n_660), .B (n_682), .C (n_548), .D (n_300), .Q
       (n_860));
  AN21X1 g50811(.A (n_681), .B (n_645), .C (n_686), .Q (n_859));
  ON22X1 g50812(.A (n_669), .B (n_685), .C (n_546), .D (n_305), .Q
       (n_858));
  AN21X1 g50813(.A (n_724), .B (n_6628), .C (n_787), .Q (n_857));
  AO22X1 g50814(.A (n_726), .B (n_641), .C (n_724), .D
       (\rs1_data[27]_39286 ), .Q (n_856));
  AN22X1 g50815(.A (n_684), .B (n_115), .C (n_124), .D (n_6628), .Q
       (n_855));
  MU2IX1 g50816(.S (n_6620), .IN0 (n_543), .IN1 (n_5542), .Q (n_854));
  ON32X1 g50817(.A (n_185), .B (n_178), .C (n_578), .D (n_639), .E
       (n_727), .Q (n_853));
  OA211X1 g50818(.A (n_642), .B (alu_2nd_operand[1]), .C (n_607), .D
       (n_627), .Q (n_883));
  AN31X1 g50819(.A (n_6458), .B (n_201), .C (n_551), .D (n_820), .Q
       (n_882));
  ON211X1 g50820(.A (n_640), .B (alu_2nd_operand[1]), .C (n_631), .D
       (n_604), .Q (n_880));
  OA211X1 g50821(.A (n_643), .B (alu_2nd_operand[1]), .C (n_608), .D
       (n_649), .Q (n_879));
  NO2X1 g50822(.A (n_792), .B (n_683), .Q (n_878));
  ON211X1 g50823(.A (n_639), .B (alu_2nd_operand[1]), .C (n_635), .D
       (n_612), .Q (n_877));
  AO222X1 g50824(.A (alu_2nd_operand[1]), .B (n_576), .C
       (\rs1_data[28]_39296 ), .D (n_127), .E (\rs1_data[29]_39336 ),
       .F (n_275), .Q (n_876));
  AN222X1 g50825(.A (n_577), .B (alu_2nd_operand[1]), .C (n_6628), .D
       (n_275), .E (n_6757), .F (n_127), .Q (n_875));
  AND2X1 g50826(.A (n_119), .B (n_6456), .Q (n_874));
  AND2X1 g50827(.A (n_119), .B (n_6458), .Q (n_872));
  NA2X1 g50830(.A (n_119), .B (n_6455), .Q (n_870));
  NA2X1 g50831(.A (n_119), .B (n_6457), .Q (n_869));
  INX1 g50832(.A (n_851), .Q (n_852));
  INX1 g50833(.A (n_848), .Q (n_849));
  INX1 g50834(.A (n_843), .Q (n_844));
  INX1 g50835(.A (n_838), .Q (n_839));
  INX1 g50836(.A (n_833), .Q (n_834));
  INX1 g50837(.A (n_830), .Q (n_831));
  INX1 g50838(.A (n_818), .Q (n_817));
  INX1 g50839(.A (n_808), .Q (n_807));
  INX1 g50840(.A (n_805), .Q (n_804));
  INX1 g50841(.A (n_800), .Q (n_801));
  OA211X1 g50842(.A (n_273), .B (n_186), .C (n_603), .D (n_630), .Q
       (n_798));
  NA2X1 g50843(.A (n_722), .B (read_data[11]), .Q (n_797));
  AO22X1 g50844(.A (n_571), .B (read_data[26]), .C (n_570), .D
       (read_data[10]), .Q (n_796));
  AN222X1 g50845(.A (n_5604), .B (n_509), .C (program_counter[0]), .D
       (n_6217), .E (n_175), .F (n_4534), .Q (n_795));
  AN222X1 g50846(.A (n_5573), .B (n_509), .C (program_counter[1]), .D
       (n_6217), .E (n_175), .F (n_6724), .Q (n_794));
  ON221X1 g50847(.A (n_183), .B (n_274), .C (n_191), .D (n_276), .E
       (n_699), .Q (n_851));
  AND4X1 g50849(.A (n_592), .B (n_652), .C (n_612), .D (n_623), .Q
       (n_850));
  AND4X1 g50850(.A (n_658), .B (n_604), .C (n_625), .D (n_616), .Q
       (n_848));
  AND4X1 g50852(.A (n_667), .B (n_591), .C (n_625), .D (n_624), .Q
       (n_846));
  AND4X1 g50853(.A (n_646), .B (n_629), .C (n_606), .D (n_619), .Q
       (n_845));
  ON211X1 g50854(.A (n_276), .B (n_194), .C (n_703), .D (n_611), .Q
       (n_843));
  AND4X1 g50855(.A (n_590), .B (n_610), .C (n_632), .D (n_677), .Q
       (n_842));
  AND4X1 g50856(.A (n_668), .B (n_598), .C (n_674), .D (n_616), .Q
       (n_841));
  AND4X1 g50857(.A (n_675), .B (n_595), .C (n_629), .D (n_659), .Q
       (n_840));
  ON211X1 g50858(.A (n_271), .B (n_186), .C (n_700), .D (n_633), .Q
       (n_838));
  ON211X1 g50859(.A (n_271), .B (n_185), .C (n_630), .D (n_701), .Q
       (n_837));
  AND4X1 g50860(.A (n_665), .B (n_589), .C (n_628), .D (n_662), .Q
       (n_836));
  ON211X1 g50861(.A (n_276), .B (n_182), .C (n_709), .D (n_603), .Q
       (n_835));
  AND4X1 g50862(.A (n_602), .B (n_592), .C (n_613), .D (n_670), .Q
       (n_833));
  NA4X1 g50863(.A (n_584), .B (n_651), .C (n_609), .D (n_664), .Q
       (n_832));
  AND4X1 g50864(.A (n_597), .B (n_585), .C (n_652), .D (n_678), .Q
       (n_830));
  AND4X1 g50865(.A (n_584), .B (n_610), .C (n_638), .D (n_676), .Q
       (n_829));
  AND4X1 g50866(.A (n_637), .B (n_607), .C (n_628), .D (n_659), .Q
       (n_828));
  AND4X1 g50867(.A (n_599), .B (n_595), .C (n_636), .D (n_617), .Q
       (n_827));
  AND4X1 g50868(.A (n_654), .B (n_626), .C (n_605), .D (n_620), .Q
       (n_826));
  AND4X1 g50869(.A (n_593), .B (n_634), .C (n_614), .D (n_621), .Q
       (n_825));
  AND4X1 g50870(.A (n_673), .B (n_601), .C (n_658), .D (n_653), .Q
       (n_824));
  AND4X1 g50871(.A (n_587), .B (n_638), .C (n_615), .D (n_679), .Q
       (n_823));
  AND4X1 g50872(.A (n_596), .B (n_588), .C (n_644), .D (n_623), .Q
       (n_822));
  OA211X1 g50873(.A (n_274), .B (n_184), .C (n_662), .D (n_698), .Q
       (n_821));
  AND3X1 g50874(.A (n_729), .B (n_201), .C (n_6459), .Q (n_820));
  NA4X1 g50875(.A (n_596), .B (n_634), .C (n_586), .D (n_666), .Q
       (n_819));
  AND4X1 g50876(.A (n_668), .B (n_636), .C (n_626), .D (n_619), .Q
       (n_818));
  AND4X1 g50877(.A (n_600), .B (n_637), .C (n_606), .D (n_656), .Q
       (n_816));
  AND4X1 g50878(.A (n_673), .B (n_598), .C (n_654), .D (n_617), .Q
       (n_815));
  AND4X1 g50879(.A (n_593), .B (n_613), .C (n_644), .D (n_622), .Q
       (n_814));
  AND4X1 g50881(.A (n_587), .B (n_608), .C (n_632), .D (n_664), .Q
       (n_812));
  NA3X1 g50882(.A (n_702), .B (n_591), .C (n_631), .Q (n_811));
  AND4X1 g50884(.A (n_599), .B (n_646), .C (n_605), .D (n_618), .Q
       (n_809));
  AND4X1 g50885(.A (n_586), .B (n_650), .C (n_609), .D (n_622), .Q
       (n_808));
  AND4X1 g50886(.A (n_594), .B (n_614), .C (n_650), .D (n_676), .Q
       (n_806));
  AND4X1 g50887(.A (n_602), .B (n_597), .C (n_588), .D (n_621), .Q
       (n_805));
  AND4X1 g50888(.A (n_594), .B (n_615), .C (n_651), .D (n_666), .Q
       (n_803));
  AND4X1 g50889(.A (n_665), .B (n_675), .C (n_600), .D (n_618), .Q
       (n_802));
  AND4X1 g50890(.A (n_667), .B (n_674), .C (n_601), .D (n_620), .Q
       (n_800));
  AO21X1 g50891(.A (n_6461), .B (n_287), .C (n_722), .Q (n_799));
  INX1 g50892(.A (n_119), .Q (n_789));
  NO2X1 g50898(.A (n_727), .B (n_647), .Q (n_787));
  ON21X1 g50899(.A (n_583), .B (n_6597), .C (n_6605), .Q (n_786));
  AN31X1 g50900(.A (n_5607), .B (n_114), .C (n_205), .D (n_6620), .Q
       (n_785));
  NO2X1 g50901(.A (n_117), .B (n_130), .Q (n_784));
  ON211X1 g50918(.A (alu_2nd_operand[1]), .B (n_285), .C (n_611), .D
       (n_633), .Q (n_783));
  OA211X1 g50936(.A (n_274), .B (n_187), .C (n_677), .D (n_690), .Q
       (n_793));
  NA3I1X1 g50938(.B (n_661), .C (n_556), .AN (n_730), .Q (n_792));
  AO222X1 g50939(.A (n_4485), .B (n_275), .C (\rs1_data[29]_39336 ), .D
       (n_127), .E (alu_2nd_operand[1]), .F (n_286), .Q (n_791));
  AN221X1 g50940(.A (alu_2nd_operand[1]), .B (n_281), .C (n_6628), .D
       (n_127), .E (n_672), .Q (n_790));
  NO2X1 g50942(.A (n_728), .B (n_6561), .Q (n_788));
  OR4X1 g50943(.A (n_5627), .B (n_6504), .C (n_6503), .D (n_6505), .Q
       (n_782));
  AN21X1 g50944(.A (n_539), .B (n_379), .C (n_123), .Q (n_781));
  AN21X1 g50945(.A (n_510), .B (n_359), .C (n_123), .Q (n_780));
  AN21X1 g50946(.A (n_533), .B (n_357), .C (n_123), .Q (n_779));
  AN21X1 g50947(.A (n_514), .B (n_376), .C (n_123), .Q (n_778));
  AN21X1 g50948(.A (n_515), .B (n_375), .C (n_123), .Q (n_777));
  AN21X1 g50949(.A (n_526), .B (n_353), .C (n_123), .Q (n_776));
  AN21X1 g50950(.A (n_528), .B (n_363), .C (n_123), .Q (n_775));
  AN21X1 g50951(.A (n_529), .B (n_362), .C (n_123), .Q (n_774));
  AN21X1 g50952(.A (n_531), .B (n_360), .C (n_123), .Q (n_773));
  AN21X1 g50953(.A (n_511), .B (n_378), .C (n_123), .Q (n_772));
  AN21X1 g50954(.A (n_516), .B (n_374), .C (n_123), .Q (n_771));
  AN21X1 g50955(.A (n_517), .B (n_373), .C (n_123), .Q (n_770));
  AN21X1 g50956(.A (n_518), .B (n_372), .C (n_123), .Q (n_769));
  AN21X1 g50957(.A (n_522), .B (n_368), .C (n_123), .Q (n_768));
  AN21X1 g50958(.A (n_523), .B (n_367), .C (n_123), .Q (n_767));
  AN21X1 g50959(.A (n_527), .B (n_364), .C (n_123), .Q (n_766));
  AN21X1 g50960(.A (n_530), .B (n_361), .C (n_123), .Q (n_765));
  AN21X1 g50961(.A (n_532), .B (n_358), .C (n_123), .Q (n_764));
  AN21X1 g50962(.A (n_534), .B (n_356), .C (n_123), .Q (n_763));
  AN21X1 g50963(.A (n_537), .B (n_354), .C (n_123), .Q (n_762));
  AN21X1 g50964(.A (n_538), .B (n_352), .C (n_123), .Q (n_761));
  AN21X1 g50965(.A (n_512), .B (n_377), .C (n_123), .Q (n_760));
  AN21X1 g50966(.A (n_513), .B (n_351), .C (n_123), .Q (n_759));
  AN21X1 g50967(.A (n_519), .B (n_371), .C (n_123), .Q (n_758));
  AN21X1 g50968(.A (n_520), .B (n_370), .C (n_123), .Q (n_757));
  AN21X1 g50969(.A (n_521), .B (n_369), .C (n_123), .Q (n_756));
  AN21X1 g50970(.A (n_524), .B (n_366), .C (n_123), .Q (n_755));
  AN21X1 g50971(.A (n_525), .B (n_365), .C (n_123), .Q (n_754));
  AN21X1 g50972(.A (n_535), .B (n_380), .C (n_123), .Q (n_753));
  AN21X1 g50973(.A (n_536), .B (n_355), .C (n_123), .Q (n_752));
  OA21X1 g50974(.A (n_350), .B (flush_37507), .C (n_122), .Q (n_751));
  NO4I2X1 g50975(.C (flush_37507), .D (n_123), .AN (n_175), .BN (mret),
       .Q (n_750));
  AN22X1 g50976(.A (n_509), .B (n_5705), .C (n_6217), .D
       (program_counter[12]), .Q (n_749));
  AN22X1 g50977(.A (n_509), .B (n_5698), .C (n_6217), .D
       (program_counter[15]), .Q (n_748));
  AN22X1 g50978(.A (n_509), .B (n_5694), .C (n_6217), .D
       (program_counter[17]), .Q (n_747));
  AN22X1 g50979(.A (n_509), .B (n_5719), .C (n_6217), .D
       (program_counter[26]), .Q (n_746));
  AN22X1 g50980(.A (n_509), .B (n_5688), .C (n_6217), .D
       (program_counter[20]), .Q (n_745));
  AN22X1 g50981(.A (n_509), .B (n_5720), .C (n_6217), .D
       (program_counter[25]), .Q (n_744));
  AN22X1 g50982(.A (n_509), .B (n_5709), .C (n_6217), .D
       (program_counter[8]), .Q (n_743));
  AN22X1 g50983(.A (n_509), .B (n_5711), .C (n_6217), .D
       (program_counter[6]), .Q (n_742));
  AN22X1 g50984(.A (n_509), .B (n_5710), .C (n_6217), .D
       (program_counter[7]), .Q (n_741));
  AN22X1 g50985(.A (n_509), .B (n_5706), .C (n_6217), .D
       (program_counter[11]), .Q (n_740));
  AN22X1 g50986(.A (n_509), .B (n_5702), .C (n_6217), .D
       (program_counter[13]), .Q (n_739));
  AN22X1 g50987(.A (n_509), .B (n_5700), .C (n_6217), .D
       (program_counter[14]), .Q (n_738));
  AN22X1 g50988(.A (n_509), .B (n_5696), .C (n_6217), .D
       (program_counter[16]), .Q (n_737));
  AN22X1 g50989(.A (n_509), .B (n_5692), .C (n_6217), .D
       (program_counter[18]), .Q (n_736));
  AN22X1 g50990(.A (n_509), .B (n_5690), .C (n_6217), .D
       (program_counter[19]), .Q (n_735));
  AN22X1 g50991(.A (n_509), .B (n_5712), .C (n_6217), .D
       (program_counter[5]), .Q (n_734));
  AN22X1 g50992(.A (n_509), .B (n_5686), .C (n_6217), .D
       (program_counter[21]), .Q (n_733));
  AN22X1 g50993(.A (n_509), .B (n_5684), .C (n_6217), .D
       (program_counter[22]), .Q (n_732));
  AN22X1 g50994(.A (n_509), .B (n_5722), .C (n_6217), .D
       (program_counter[23]), .Q (n_731));
  INX1 g50996(.A (n_727), .Q (n_726));
  AN22X1 g50997(.A (n_509), .B (n_5721), .C (n_6217), .D
       (program_counter[24]), .Q (n_721));
  AN22X1 g50998(.A (n_509), .B (n_5717), .C (n_6217), .D
       (program_counter[28]), .Q (n_720));
  AN22X1 g50999(.A (n_509), .B (n_5718), .C (n_6217), .D
       (program_counter[27]), .Q (n_719));
  AN22X1 g51000(.A (n_509), .B (n_5715), .C (n_6217), .D
       (program_counter[29]), .Q (n_718));
  AN22X1 g51001(.A (n_509), .B (n_5716), .C (n_6217), .D
       (program_counter[2]), .Q (n_717));
  AN22X1 g51002(.A (n_509), .B (n_5704), .C (n_6217), .D
       (program_counter[30]), .Q (n_716));
  AN22X1 g51003(.A (n_509), .B (n_5682), .C (n_6217), .D
       (program_counter[31]), .Q (n_715));
  AN22X1 g51004(.A (n_509), .B (n_5714), .C (n_6217), .D
       (program_counter[3]), .Q (n_714));
  AN22X1 g51005(.A (n_509), .B (n_5708), .C (n_6217), .D
       (program_counter[9]), .Q (n_713));
  AN22X1 g51006(.A (n_509), .B (n_5713), .C (n_6217), .D
       (program_counter[4]), .Q (n_712));
  AN22X1 g51007(.A (n_509), .B (n_5707), .C (n_6217), .D
       (program_counter[10]), .Q (n_711));
  NO2X1 g51009(.A (n_562), .B (n_123), .Q (n_710));
  OA21X1 g51010(.A (n_274), .B (n_199), .C (n_624), .Q (n_709));
  ON32X1 g51014(.A (n_190), .B (alu_2nd_operand[8]), .C (n_297), .D
       (n_200), .E (alu_2nd_operand[9]), .Q (n_705));
  AN221X1 g51015(.A (n_190), .B (alu_2nd_operand[8]), .C
       (alu_2nd_operand[7]), .D (n_196), .E (n_297), .Q (n_704));
  OA21X1 g51016(.A (n_274), .B (n_182), .C (n_678), .Q (n_703));
  OA21X1 g51017(.A (n_271), .B (n_199), .C (n_653), .Q (n_702));
  AN22X1 g51018(.A (n_127), .B (\rs1_data[26]_39276 ), .C (n_275), .D
       (\rs1_data[27]_39286 ), .Q (n_701));
  AN22X1 g51019(.A (n_127), .B (\rs1_data[27]_39286 ), .C (n_275), .D
       (\rs1_data[28]_39296 ), .Q (n_700));
  AN22X1 g51020(.A (n_127), .B (n_4461), .C (n_272), .D (n_6628), .Q
       (n_699));
  AN22X1 g51021(.A (n_128), .B (n_4465), .C (n_272), .D (n_6757), .Q
       (n_698));
  AN22X1 g51022(.A (n_128), .B (n_6628), .C (n_272), .D (n_6629), .Q
       (n_697));
  NO2X1 g51023(.A (n_550), .B (n_123), .Q (n_696));
  NO2X1 g51024(.A (n_560), .B (n_123), .Q (n_695));
  NO2X1 g51025(.A (n_541), .B (n_123), .Q (n_694));
  NO2X1 g51026(.A (n_540), .B (n_123), .Q (n_693));
  NO2X1 g51027(.A (n_542), .B (n_123), .Q (n_692));
  NA2X1 g51028(.A (n_581), .B (n_281), .Q (n_691));
  AN22X1 g51029(.A (n_128), .B (n_4461), .C (n_272), .D (n_4465), .Q
       (n_690));
  ON32X1 g51030(.A (n_189), .B (alu_2nd_operand[24]), .C (n_312), .D
       (n_199), .E (alu_2nd_operand[25]), .Q (n_689));
  NO3I1X1 g51031(.B (n_669), .C (n_309), .AN (n_340), .Q (n_688));
  AN21X1 g51032(.A (n_281), .B (n_179), .C (n_672), .Q (n_687));
  AN21X1 g51033(.A (n_317), .B (n_331), .C (n_295), .Q (n_686));
  AN31X1 g51034(.A (n_4484), .B (n_207), .C (n_308), .D (n_318), .Q
       (n_685));
  ON21X1 g51035(.A (n_335), .B (n_329), .C (n_293), .Q (n_684));
  NA3X1 g51036(.A (n_645), .B (n_116), .C (n_314), .Q (n_683));
  ON31X1 g51037(.A (n_181), .B (alu_2nd_operand[28]), .C (n_301), .D
       (n_321), .Q (n_682));
  ON21X1 g51038(.A (n_320), .B (n_313), .C (n_341), .Q (n_681));
  ON211X1 g51039(.A (n_209), .B (\rs1_data[28]_39296 ), .C (n_302), .D
       (n_660), .Q (n_730));
  ON221X1 g51040(.A (n_174), .B (n_6065), .C (n_173), .D (n_6064), .E
       (n_565), .Q (n_729));
  OR4X1 g51041(.A (jalr_type), .B (n_201), .C (jal_type), .D (n_270),
       .Q (n_728));
  NA2X1 g51042(.A (n_573), .B (alu_2nd_operand[1]), .Q (n_727));
  NO2X1 g51044(.A (n_578), .B (n_4533), .Q (n_724));
  OR2X1 g51045(.A (n_563), .B (n_569), .Q (n_723));
  NO2X1 g51046(.A (n_561), .B (n_6367), .Q (n_722));
  INX1 g51053(.A (n_640), .Q (n_641));
  INX1 g51054(.A (n_575), .Q (n_574));
  INX1 g51055(.A (n_573), .Q (n_572));
  INX1 g51057(.A (n_129), .Q (n_568));
  NA2X1 g51059(.A (n_5707), .B (n_270), .Q (n_567));
  NA2X1 g51060(.A (n_5706), .B (n_270), .Q (n_566));
  AN22X1 g51061(.A (n_212), .B (read_data[15]), .C (n_6461), .D
       (read_data[7]), .Q (n_565));
  NO3X1 g51062(.A (n_175), .B (flush_37507), .C (n_123), .Q (n_564));
  NO2I1X1 g51063(.B (n_6065), .AN (n_287), .Q (n_563));
  MU2IX1 g51065(.S (n_6373), .IN0 (csr_mcause_code[2]), .IN1 (n_5988),
       .Q (n_562));
  AN21X1 g51088(.A (n_204), .B (n_5606), .C (n_6721), .Q (n_561));
  MU2IX1 g51097(.S (n_6373), .IN0 (csr_mcause_code[4]), .IN1 (n_4535),
       .Q (n_560));
  AN21X1 g51129(.A (n_5607), .B (n_6373), .C (n_6071), .Q (n_559));
  NO2I1X1 g51130(.B (n_295), .AN (n_331), .Q (n_558));
  AND2X1 g51131(.A (n_317), .B (n_316), .Q (n_557));
  AN21X1 g51132(.A (alu_2nd_operand[24]), .B (n_189), .C (n_312), .Q
       (n_556));
  NO2X1 g51133(.A (n_318), .B (n_309), .Q (n_555));
  ON22X1 g51134(.A (alu_2nd_operand[11]), .B (n_202), .C
       (alu_2nd_operand[10]), .D (n_195), .Q (n_554));
  ON22X1 g51135(.A (alu_2nd_operand[27]), .B (n_194), .C
       (alu_2nd_operand[26]), .D (n_182), .Q (n_553));
  AND2X1 g51136(.A (n_320), .B (n_116), .Q (n_552));
  MU2X1 g51137(.S (n_5573), .IN0 (read_data[15]), .IN1 (read_data[31]),
       .Q (n_551));
  MU2IX1 g51138(.S (n_6373), .IN0 (csr_mcause_code[1]), .IN1 (n_6724),
       .Q (n_550));
  AND2X1 g51139(.A (n_341), .B (n_314), .Q (n_549));
  ON21X1 g51140(.A (alu_2nd_operand[30]), .B (n_186), .C (n_322), .Q
       (n_548));
  NO2X1 g51141(.A (n_323), .B (n_330), .Q (n_547));
  NO2X1 g51142(.A (n_332), .B (n_323), .Q (n_546));
  AND2X1 g51143(.A (n_321), .B (n_302), .Q (n_545));
  NO2X1 g51144(.A (n_332), .B (n_305), .Q (n_544));
  AO21X1 g51145(.A (n_211), .B (n_4549), .C (n_5987), .Q (n_543));
  MU2IX1 g51146(.S (n_6373), .IN0 (csr_mcause_code[3]), .IN1 (n_5987),
       .Q (n_542));
  MU2IX1 g51147(.S (n_6373), .IN0 (csr_mcause_interrupt_flag), .IN1
       (n_5985), .Q (n_541));
  MU2IX1 g51148(.S (n_6373), .IN0 (csr_mcause_code[0]), .IN1 (n_4534),
       .Q (n_540));
  NA2X1 g51149(.A (n_127), .B (n_4487), .Q (n_679));
  NA2X1 g51150(.A (n_127), .B (n_4481), .Q (n_678));
  NA2X1 g51151(.A (n_127), .B (n_4460), .Q (n_677));
  NA2X1 g51152(.A (n_127), .B (n_4476), .Q (n_676));
  NA2X1 g51153(.A (n_275), .B (n_4474), .Q (n_675));
  NA2X1 g51154(.A (n_275), .B (n_4477), .Q (n_674));
  NA2X1 g51155(.A (n_272), .B (n_4477), .Q (n_673));
  NO2X1 g51156(.A (n_293), .B (n_4533), .Q (n_672));
  NA2X1 g51157(.A (n_127), .B (\rs1_data[23]_39246 ), .Q (n_670));
  OR2X1 g51158(.A (n_305), .B (n_330), .Q (n_669));
  NA2X1 g51159(.A (n_272), .B (n_4482), .Q (n_668));
  NA2X1 g51160(.A (n_272), .B (n_4479), .Q (n_667));
  NA2X1 g51161(.A (n_127), .B (\rs1_data[15]_39476 ), .Q (n_666));
  NA2X1 g51162(.A (n_272), .B (n_4487), .Q (n_665));
  NA2X1 g51163(.A (n_127), .B (n_4474), .Q (n_664));
  AN21X1 g51164(.A (alu_2nd_operand[10]), .B (n_195), .C (n_306), .Q
       (n_663));
  NA2X1 g51165(.A (n_127), .B (n_4466), .Q (n_662));
  AN21X1 g51166(.A (alu_2nd_operand[26]), .B (n_182), .C (n_303), .Q
       (n_661));
  AN21X1 g51167(.A (alu_2nd_operand[30]), .B (n_186), .C (n_299), .Q
       (n_660));
  NA2X1 g51168(.A (n_127), .B (n_4480), .Q (n_659));
  NA2X1 g51169(.A (n_275), .B (n_4479), .Q (n_658));
  NA2X1 g51170(.A (n_127), .B (n_4464), .Q (n_656));
  NA2X1 g51171(.A (n_278), .B (alu_2nd_operand[4]), .Q (n_655));
  NA2X1 g51172(.A (n_275), .B (n_4482), .Q (n_654));
  NA2X1 g51173(.A (n_127), .B (n_4463), .Q (n_653));
  NA2X1 g51174(.A (n_128), .B (\rs1_data[23]_39246 ), .Q (n_652));
  NA2X1 g51175(.A (n_128), .B (n_4476), .Q (n_651));
  NA2X1 g51176(.A (n_128), .B (\rs1_data[15]_39476 ), .Q (n_650));
  NA2X1 g51177(.A (n_128), .B (n_4460), .Q (n_649));
  MU2IX1 g51178(.S (n_4533), .IN0 (n_6757), .IN1 (n_6628), .Q (n_648));
  MU2IX1 g51179(.S (n_4533), .IN0 (n_4465), .IN1 (n_6757), .Q (n_647));
  NA2X1 g51180(.A (n_275), .B (n_4476), .Q (n_646));
  NO2X1 g51181(.A (n_315), .B (n_295), .Q (n_645));
  NA2X1 g51182(.A (n_128), .B (n_4477), .Q (n_644));
  MU2IX1 g51183(.S (n_4533), .IN0 (n_4466), .IN1 (n_4461), .Q (n_643));
  MU2IX1 g51184(.S (n_4533), .IN0 (n_4461), .IN1 (n_4465), .Q (n_642));
  MU2IX1 g51185(.S (n_4533), .IN0 (n_4481), .IN1 (\rs1_data[26]_39276
       ), .Q (n_640));
  MU2IX1 g51186(.S (n_4533), .IN0 (\rs1_data[26]_39276 ), .IN1
       (\rs1_data[27]_39286 ), .Q (n_639));
  NA2X1 g51187(.A (n_128), .B (n_4474), .Q (n_638));
  NA2X1 g51188(.A (n_275), .B (n_4487), .Q (n_637));
  NA2X1 g51189(.A (n_275), .B (\rs1_data[15]_39476 ), .Q (n_636));
  NA2X1 g51190(.A (n_128), .B (n_4481), .Q (n_635));
  NA2X1 g51191(.A (n_128), .B (n_4482), .Q (n_634));
  NA2X1 g51192(.A (n_128), .B (\rs1_data[29]_39336 ), .Q (n_633));
  NA2X1 g51193(.A (n_128), .B (n_4487), .Q (n_632));
  NA2X1 g51194(.A (n_128), .B (n_4483), .Q (n_631));
  NA2X1 g51195(.A (n_128), .B (\rs1_data[28]_39296 ), .Q (n_630));
  NA2X1 g51196(.A (n_128), .B (n_4475), .Q (n_629));
  NA2X1 g51197(.A (n_128), .B (n_4464), .Q (n_628));
  NA2X1 g51198(.A (n_128), .B (n_4466), .Q (n_627));
  NA2X1 g51199(.A (n_128), .B (n_4484), .Q (n_626));
  NA2X1 g51200(.A (n_128), .B (n_4463), .Q (n_625));
  NA2X1 g51201(.A (n_127), .B (n_4483), .Q (n_624));
  NA2X1 g51202(.A (n_127), .B (n_4479), .Q (n_623));
  NA2X1 g51203(.A (n_127), .B (n_4482), .Q (n_622));
  NA2X1 g51204(.A (n_127), .B (n_4477), .Q (n_621));
  NA2X1 g51205(.A (n_127), .B (n_4478), .Q (n_620));
  NA2X1 g51206(.A (n_127), .B (\rs1_data[14]_39466 ), .Q (n_619));
  NA2X1 g51207(.A (n_127), .B (n_4475), .Q (n_618));
  NA2X1 g51208(.A (n_127), .B (n_4484), .Q (n_617));
  NA2X1 g51209(.A (n_127), .B (n_4486), .Q (n_616));
  NA2X1 g51210(.A (n_272), .B (n_4475), .Q (n_615));
  NA2X1 g51211(.A (n_272), .B (n_4484), .Q (n_614));
  NA2X1 g51212(.A (n_272), .B (n_4486), .Q (n_613));
  NA2X1 g51213(.A (n_272), .B (n_4483), .Q (n_612));
  NA2X1 g51214(.A (n_272), .B (\rs1_data[28]_39296 ), .Q (n_611));
  NA2X1 g51215(.A (n_272), .B (n_4480), .Q (n_610));
  NA2X1 g51216(.A (n_272), .B (\rs1_data[14]_39466 ), .Q (n_609));
  NA2X1 g51217(.A (n_272), .B (n_4464), .Q (n_608));
  NA2X1 g51218(.A (n_272), .B (n_4460), .Q (n_607));
  NA2X1 g51219(.A (n_272), .B (n_4474), .Q (n_606));
  NA2X1 g51220(.A (n_272), .B (\rs1_data[15]_39476 ), .Q (n_605));
  NA2X1 g51221(.A (n_272), .B (\rs1_data[23]_39246 ), .Q (n_604));
  NA2X1 g51222(.A (n_272), .B (\rs1_data[27]_39286 ), .Q (n_603));
  NA2X1 g51223(.A (n_128), .B (n_4479), .Q (n_602));
  NA2X1 g51224(.A (n_128), .B (n_4486), .Q (n_601));
  NA2X1 g51225(.A (n_128), .B (n_4480), .Q (n_600));
  NA2X1 g51226(.A (n_128), .B (\rs1_data[14]_39466 ), .Q (n_599));
  NA2X1 g51227(.A (n_128), .B (n_4478), .Q (n_598));
  NA2X1 g51228(.A (n_272), .B (n_4463), .Q (n_597));
  NA2X1 g51229(.A (n_272), .B (n_4478), .Q (n_596));
  NA2X1 g51230(.A (n_272), .B (n_4476), .Q (n_595));
  NA2X1 g51231(.A (n_275), .B (\rs1_data[14]_39466 ), .Q (n_594));
  NA2X1 g51232(.A (n_275), .B (n_4478), .Q (n_593));
  NA2X1 g51233(.A (n_275), .B (n_4463), .Q (n_592));
  NA2X1 g51234(.A (n_275), .B (\rs1_data[23]_39246 ), .Q (n_591));
  NA2X1 g51235(.A (n_275), .B (n_4464), .Q (n_590));
  NA2X1 g51236(.A (n_275), .B (n_4460), .Q (n_589));
  NA2X1 g51237(.A (n_275), .B (n_4486), .Q (n_588));
  NA2X1 g51238(.A (n_275), .B (n_4480), .Q (n_587));
  NA2X1 g51239(.A (n_275), .B (n_4484), .Q (n_586));
  NA2X1 g51240(.A (n_275), .B (n_4483), .Q (n_585));
  NA2X1 g51241(.A (n_275), .B (n_4475), .Q (n_584));
  NA2X1 g51242(.A (n_322), .B (n_300), .Q (n_583));
  AND2X1 g51249(.A (n_288), .B (alu_2nd_operand[3]), .Q (n_582));
  AND2X1 g51250(.A (n_288), .B (n_294), .Q (n_581));
  NA2X1 g51251(.A (n_282), .B (n_124), .Q (n_580));
  NA2X1 g51252(.A (n_282), .B (alu_2nd_operand[2]), .Q (n_579));
  NA2X1 g51253(.A (n_288), .B (n_310), .Q (n_578));
  AO21X1 g51254(.A (n_4533), .B (n_6629), .C (n_333), .Q (n_577));
  MU2IX1 g51255(.S (n_4533), .IN0 (n_198), .IN1 (n_186), .Q (n_576));
  AND2X1 g51256(.A (n_283), .B (n_180), .Q (n_575));
  NO2X1 g51257(.A (n_279), .B (alu_2nd_operand[4]), .Q (n_573));
  NO2I1X1 g51258(.B (n_6064), .AN (n_287), .Q (n_571));
  NO2I1X1 g51259(.B (n_6067), .AN (n_287), .Q (n_570));
  AND3X1 g51260(.A (n_5573), .B (n_201), .C (n_5606), .Q (n_569));
  AND2X1 g51469(.A (rw_address[28]), .B (n_122), .Q (n_508));
  AND2X1 g51470(.A (rw_address[16]), .B (n_121), .Q (n_507));
  AND2X1 g51471(.A (rw_address[12]), .B (n_121), .Q (n_506));
  AND2X1 g51472(.A (rw_address[25]), .B (n_122), .Q (n_505));
  AND2X1 g51473(.A (rw_address[13]), .B (n_121), .Q (n_504));
  AND2X1 g51474(.A (rw_address[14]), .B (n_122), .Q (n_503));
  AND2X1 g51475(.A (rw_address[11]), .B (n_122), .Q (n_502));
  AND2X1 g51476(.A (rw_address[15]), .B (n_122), .Q (n_501));
  AND2X1 g51477(.A (rw_address[5]), .B (n_121), .Q (n_500));
  AND2X1 g51478(.A (rw_address[10]), .B (n_121), .Q (n_499));
  AND2X1 g51479(.A (rw_address[26]), .B (n_122), .Q (n_498));
  AND2X1 g51480(.A (rw_address[9]), .B (n_122), .Q (n_497));
  AND2X1 g51481(.A (rw_address[8]), .B (n_121), .Q (n_496));
  AND2X1 g51482(.A (rw_address[1]), .B (n_121), .Q (n_495));
  AND2X1 g51483(.A (rw_address[21]), .B (n_121), .Q (n_494));
  AND2X1 g51484(.A (rw_address[18]), .B (n_122), .Q (n_493));
  AND2X1 g51485(.A (rw_address[22]), .B (n_122), .Q (n_492));
  AND2X1 g51486(.A (rw_address[29]), .B (n_122), .Q (n_491));
  AND2X1 g51487(.A (rw_address[27]), .B (n_121), .Q (n_490));
  AND2X1 g51488(.A (rw_address[23]), .B (n_121), .Q (n_489));
  AND2X1 g51489(.A (rw_address[24]), .B (n_121), .Q (n_488));
  AND2X1 g51490(.A (rw_address[20]), .B (n_121), .Q (n_487));
  AND2X1 g51491(.A (rw_address[17]), .B (n_121), .Q (n_486));
  AND2X1 g51492(.A (rw_address[19]), .B (n_122), .Q (n_485));
  AND2X1 g51493(.A (rw_address[31]), .B (n_122), .Q (n_484));
  AND2X1 g51494(.A (rw_address[30]), .B (n_121), .Q (n_483));
  AND2X1 g51495(.A (rw_address[4]), .B (n_121), .Q (n_482));
  AND2X1 g51496(.A (rw_address[2]), .B (n_122), .Q (n_481));
  AND2X1 g51497(.A (rw_address[6]), .B (n_121), .Q (n_480));
  AND2X1 g51498(.A (rw_address[3]), .B (n_122), .Q (n_479));
  AND2X1 g51499(.A (rw_address[7]), .B (n_121), .Q (n_478));
  AND2X1 g51500(.A (rw_address[0]), .B (n_121), .Q (n_477));
  AND2X1 g51501(.A (write_strobe[0]), .B (n_122), .Q (n_476));
  AND2X1 g51502(.A (write_strobe[2]), .B (n_122), .Q (n_475));
  AND2X1 g51503(.A (write_strobe[1]), .B (n_122), .Q (n_474));
  AND2X1 g51504(.A (write_strobe[3]), .B (n_122), .Q (n_473));
  AND2X1 g51505(.A (instruction_address[2]), .B (n_121), .Q (n_472));
  AND2X1 g51506(.A (instruction_address[4]), .B (n_122), .Q (n_471));
  AND2X1 g51507(.A (instruction_address[3]), .B (n_122), .Q (n_470));
  AND2X1 g51508(.A (instruction_address[7]), .B (n_122), .Q (n_469));
  AND2X1 g51509(.A (instruction_address[6]), .B (n_122), .Q (n_468));
  AND2X1 g51510(.A (instruction_address[12]), .B (n_122), .Q (n_467));
  AND2X1 g51511(.A (instruction_address[14]), .B (n_122), .Q (n_466));
  AND2X1 g51512(.A (instruction_address[26]), .B (n_122), .Q (n_465));
  AND2X1 g51513(.A (instruction_address[25]), .B (n_122), .Q (n_464));
  AND2X1 g51514(.A (instruction_address[16]), .B (n_121), .Q (n_463));
  AND2X1 g51515(.A (instruction_address[9]), .B (n_121), .Q (n_462));
  AND2X1 g51516(.A (instruction_address[5]), .B (n_122), .Q (n_461));
  AND2X1 g51517(.A (instruction_address[27]), .B (n_121), .Q (n_460));
  AND2X1 g51518(.A (instruction_address[8]), .B (n_122), .Q (n_459));
  AND2X1 g51519(.A (instruction_address[13]), .B (n_122), .Q (n_458));
  AND2X1 g51520(.A (instruction_address[15]), .B (n_122), .Q (n_457));
  AND2X1 g51521(.A (instruction_address[28]), .B (n_122), .Q (n_456));
  AND2X1 g51522(.A (instruction_address[11]), .B (n_121), .Q (n_455));
  AND2X1 g51523(.A (instruction_address[10]), .B (n_121), .Q (n_454));
  AND2X1 g51524(.A (instruction_address[18]), .B (n_121), .Q (n_453));
  AND2X1 g51525(.A (instruction_address[30]), .B (n_121), .Q (n_452));
  AND2X1 g51526(.A (instruction_address[23]), .B (n_122), .Q (n_451));
  AND2X1 g51527(.A (instruction_address[19]), .B (n_122), .Q (n_450));
  AND2X1 g51528(.A (instruction_address[29]), .B (n_122), .Q (n_449));
  AND2X1 g51529(.A (instruction_address[31]), .B (n_121), .Q (n_448));
  AND2X1 g51530(.A (instruction_address[24]), .B (n_121), .Q (n_447));
  AND2X1 g51531(.A (instruction_address[22]), .B (n_121), .Q (n_446));
  AND2X1 g51532(.A (instruction_address[20]), .B (n_121), .Q (n_445));
  AND2X1 g51533(.A (instruction_address[21]), .B (n_122), .Q (n_444));
  AND2X1 g51534(.A (instruction_address[17]), .B (n_122), .Q (n_443));
  AND2X1 g51535(.A (instruction_address[1]), .B (n_121), .Q (n_442));
  AND2X1 g51536(.A (instruction_address[0]), .B (n_121), .Q (n_441));
  AND2X1 g51537(.A (write_request), .B (n_122), .Q (n_440));
  AND2X1 g51538(.A (read_request), .B (n_122), .Q (n_439));
  AND2X1 g51539(.A (n_6529), .B (n_122), .Q (n_438));
  AND2X1 g51540(.A (n_6536), .B (n_122), .Q (n_437));
  AND2X1 g51541(.A (n_6535), .B (n_122), .Q (n_436));
  AND2X1 g51542(.A (n_6533), .B (n_122), .Q (n_435));
  AND2X1 g51543(.A (n_6530), .B (n_122), .Q (n_434));
  AND2X1 g51544(.A (n_6532), .B (n_122), .Q (n_433));
  AND2X1 g51545(.A (n_6528), .B (n_122), .Q (n_432));
  AND2X1 g51546(.A (n_6526), .B (n_122), .Q (n_431));
  AND2X1 g51547(.A (n_6537), .B (n_122), .Q (n_430));
  AND2X1 g51548(.A (n_6543), .B (n_122), .Q (n_429));
  AND2X1 g51549(.A (n_6527), .B (n_122), .Q (n_428));
  AND2X1 g51550(.A (n_6540), .B (n_122), .Q (n_427));
  AND2X1 g51551(.A (n_6538), .B (n_122), .Q (n_426));
  AND2X1 g51552(.A (n_6534), .B (n_122), .Q (n_425));
  AND2X1 g51553(.A (n_6525), .B (n_122), .Q (n_424));
  AND2X1 g51554(.A (n_6539), .B (n_122), .Q (n_423));
  AND2X1 g51555(.A (n_6545), .B (n_122), .Q (n_422));
  AND2X1 g51556(.A (n_6546), .B (n_122), .Q (n_421));
  AND2X1 g51557(.A (n_6544), .B (n_122), .Q (n_420));
  AND2X1 g51558(.A (n_6524), .B (n_122), .Q (n_419));
  AND2X1 g51559(.A (n_6541), .B (n_122), .Q (n_418));
  AND2X1 g51560(.A (n_6552), .B (n_122), .Q (n_417));
  AND2X1 g51561(.A (n_6549), .B (n_122), .Q (n_416));
  AND2X1 g51562(.A (n_6522), .B (n_122), .Q (n_415));
  AND2X1 g51563(.A (n_6550), .B (n_122), .Q (n_414));
  AND2X1 g51564(.A (n_6548), .B (n_122), .Q (n_413));
  AND2X1 g51565(.A (n_6551), .B (n_122), .Q (n_412));
  AND2X1 g51566(.A (n_6553), .B (n_122), .Q (n_411));
  AND2X1 g51567(.A (n_6542), .B (n_122), .Q (n_410));
  AND2X1 g51568(.A (n_6531), .B (n_122), .Q (n_409));
  AND2X1 g51569(.A (n_6547), .B (n_122), .Q (n_408));
  AND2X1 g51570(.A (n_6523), .B (n_122), .Q (n_407));
  AND2X1 g51571(.A (n_6724), .B (n_122), .Q (n_406));
  AND2X1 g51576(.A (write_data[31]), .B (n_122), .Q (n_405));
  AND2X1 g51577(.A (write_data[30]), .B (n_121), .Q (n_404));
  AND2X1 g51578(.A (write_data[24]), .B (n_121), .Q (n_403));
  AND2X1 g51579(.A (write_data[28]), .B (n_121), .Q (n_402));
  AND2X1 g51580(.A (write_data[29]), .B (n_121), .Q (n_401));
  AND2X1 g51581(.A (write_data[25]), .B (n_121), .Q (n_400));
  AND2X1 g51582(.A (write_data[26]), .B (n_121), .Q (n_399));
  AND2X1 g51583(.A (write_data[27]), .B (n_121), .Q (n_398));
  AND2X1 g51584(.A (write_data[19]), .B (n_122), .Q (n_397));
  AND2X1 g51585(.A (write_data[23]), .B (n_122), .Q (n_396));
  AND2X1 g51586(.A (write_data[18]), .B (n_121), .Q (n_395));
  AND2X1 g51587(.A (write_data[16]), .B (n_121), .Q (n_394));
  AND2X1 g51588(.A (write_data[22]), .B (n_122), .Q (n_393));
  AND2X1 g51589(.A (write_data[21]), .B (n_122), .Q (n_392));
  AND2X1 g51590(.A (write_data[20]), .B (n_122), .Q (n_391));
  AND2X1 g51591(.A (write_data[17]), .B (n_122), .Q (n_390));
  AND2X1 g51592(.A (write_data[12]), .B (n_122), .Q (n_389));
  AND2X1 g51593(.A (write_data[8]), .B (n_122), .Q (n_388));
  AND2X1 g51594(.A (write_data[9]), .B (n_122), .Q (n_387));
  AND2X1 g51595(.A (write_data[13]), .B (n_122), .Q (n_386));
  AND2X1 g51596(.A (write_data[14]), .B (n_122), .Q (n_385));
  AND2X1 g51597(.A (write_data[10]), .B (n_121), .Q (n_384));
  AND2X1 g51598(.A (write_data[15]), .B (n_121), .Q (n_383));
  AND2X1 g51599(.A (write_data[11]), .B (n_121), .Q (n_382));
  AND2X1 g51600(.A (write_data[1]), .B (n_122), .Q (n_381));
  NA2X1 g51601(.A (take_trap_39145), .B (program_counter[6]), .Q
       (n_380));
  NA2X1 g51602(.A (take_trap_39145), .B (program_counter[10]), .Q
       (n_379));
  NA2X1 g51603(.A (take_trap_39145), .B (program_counter[11]), .Q
       (n_378));
  NA2X1 g51604(.A (take_trap_39145), .B (program_counter[12]), .Q
       (n_377));
  NA2X1 g51605(.A (take_trap_39145), .B (program_counter[14]), .Q
       (n_376));
  NA2X1 g51606(.A (take_trap_39145), .B (program_counter[15]), .Q
       (n_375));
  NA2X1 g51607(.A (take_trap_39145), .B (program_counter[16]), .Q
       (n_374));
  NA2X1 g51608(.A (take_trap_39145), .B (program_counter[17]), .Q
       (n_373));
  NA2X1 g51609(.A (take_trap_39145), .B (program_counter[18]), .Q
       (n_372));
  NA2X1 g51610(.A (take_trap_39145), .B (program_counter[19]), .Q
       (n_371));
  NA2X1 g51611(.A (take_trap_39145), .B (program_counter[20]), .Q
       (n_370));
  NA2X1 g51612(.A (take_trap_39145), .B (program_counter[21]), .Q
       (n_369));
  NA2X1 g51613(.A (take_trap_39145), .B (program_counter[22]), .Q
       (n_368));
  NA2X1 g51614(.A (take_trap_39145), .B (program_counter[23]), .Q
       (n_367));
  NA2X1 g51615(.A (take_trap_39145), .B (program_counter[24]), .Q
       (n_366));
  NA2X1 g51616(.A (take_trap_39145), .B (program_counter[25]), .Q
       (n_365));
  NA2X1 g51617(.A (take_trap_39145), .B (program_counter[27]), .Q
       (n_364));
  NA2X1 g51618(.A (take_trap_39145), .B (program_counter[28]), .Q
       (n_363));
  NA2X1 g51619(.A (take_trap_39145), .B (program_counter[29]), .Q
       (n_362));
  NA2X1 g51620(.A (take_trap_39145), .B (program_counter[2]), .Q
       (n_361));
  NA2X1 g51621(.A (take_trap_39145), .B (program_counter[30]), .Q
       (n_360));
  NA2X1 g51622(.A (take_trap_39145), .B (program_counter[31]), .Q
       (n_359));
  NA2X1 g51623(.A (take_trap_39145), .B (program_counter[3]), .Q
       (n_358));
  NA2X1 g51624(.A (take_trap_39145), .B (program_counter[4]), .Q
       (n_357));
  NA2X1 g51625(.A (take_trap_39145), .B (program_counter[5]), .Q
       (n_356));
  NA2X1 g51626(.A (take_trap_39145), .B (program_counter[7]), .Q
       (n_355));
  NA2X1 g51627(.A (take_trap_39145), .B (program_counter[9]), .Q
       (n_354));
  NA2X1 g51628(.A (take_trap_39145), .B (program_counter[26]), .Q
       (n_353));
  NA2X1 g51629(.A (take_trap_39145), .B (program_counter[8]), .Q
       (n_352));
  NA2X1 g51630(.A (take_trap_39145), .B (program_counter[13]), .Q
       (n_351));
  NO2X1 g51631(.A (take_trap_39145), .B (mret), .Q (n_350));
  NO2X1 g51632(.A (load_request_BAR), .B (n_123), .Q (n_349));
  AND2X1 g51633(.A (write_data[4]), .B (n_122), .Q (n_348));
  AND2X1 g51634(.A (write_data[7]), .B (n_121), .Q (n_347));
  AND2X1 g51635(.A (write_data[3]), .B (n_121), .Q (n_346));
  AND2X1 g51636(.A (write_data[6]), .B (n_121), .Q (n_345));
  AND2X1 g51637(.A (write_data[5]), .B (n_121), .Q (n_344));
  AND2X1 g51638(.A (write_data[0]), .B (n_122), .Q (n_343));
  AND2X1 g51639(.A (write_data[2]), .B (n_121), .Q (n_342));
  NA2X1 g51640(.A (n_175), .B (n_5749), .Q (n_539));
  NA2X1 g51641(.A (n_175), .B (n_5751), .Q (n_538));
  NA2X1 g51642(.A (n_175), .B (n_5750), .Q (n_537));
  NA2X1 g51643(.A (n_175), .B (n_6726), .Q (n_536));
  NA2X1 g51644(.A (n_175), .B (n_6730), .Q (n_535));
  NA2X1 g51645(.A (n_175), .B (n_6731), .Q (n_534));
  NA2X1 g51646(.A (n_175), .B (n_4535), .Q (n_533));
  NA2X1 g51647(.A (n_175), .B (n_5987), .Q (n_532));
  NA2X1 g51648(.A (n_175), .B (n_5729), .Q (n_531));
  NA2X1 g51649(.A (n_175), .B (n_5988), .Q (n_530));
  NA2X1 g51650(.A (n_175), .B (n_5730), .Q (n_529));
  NA2X1 g51651(.A (n_175), .B (n_5731), .Q (n_528));
  NA2X1 g51652(.A (n_175), .B (n_5732), .Q (n_527));
  NA2X1 g51653(.A (n_175), .B (n_5733), .Q (n_526));
  NA2X1 g51654(.A (n_175), .B (n_5734), .Q (n_525));
  NA2X1 g51655(.A (n_175), .B (n_5735), .Q (n_524));
  NA2X1 g51656(.A (n_175), .B (n_5736), .Q (n_523));
  NA2X1 g51657(.A (n_175), .B (n_5737), .Q (n_522));
  NA2X1 g51658(.A (n_175), .B (n_5738), .Q (n_521));
  NA2X1 g51659(.A (n_175), .B (n_5739), .Q (n_520));
  NA2X1 g51660(.A (n_175), .B (n_5740), .Q (n_519));
  NA2X1 g51661(.A (n_175), .B (n_5741), .Q (n_518));
  NA2X1 g51662(.A (n_175), .B (n_5742), .Q (n_517));
  NA2X1 g51663(.A (n_175), .B (n_5743), .Q (n_516));
  NA2X1 g51664(.A (n_175), .B (n_4538), .Q (n_515));
  NA2X1 g51665(.A (n_175), .B (n_4536), .Q (n_514));
  NA2X1 g51666(.A (n_175), .B (n_5746), .Q (n_513));
  NA2X1 g51667(.A (n_175), .B (n_5747), .Q (n_512));
  NA2X1 g51668(.A (n_175), .B (n_5748), .Q (n_511));
  NA2X1 g51669(.A (n_175), .B (n_5985), .Q (n_510));
  OR2X1 g51670(.A (n_6218), .B (n_6595), .Q (n_509));
  INX1 g51671(.A (n_336), .Q (n_337));
  INX1 g51672(.A (n_334), .Q (n_335));
  INX1 g51673(.A (n_315), .Q (n_316));
  INX1 g51674(.A (n_313), .Q (n_314));
  INX1 g51675(.A (n_311), .Q (n_312));
  INX1 g51676(.A (n_309), .Q (n_308));
  INX1 g51677(.A (n_307), .Q (n_306));
  INX1 g51678(.A (n_304), .Q (n_303));
  INX1 g51679(.A (n_302), .Q (n_301));
  INX1 g51680(.A (n_300), .Q (n_299));
  INX1 g51681(.A (n_296), .Q (n_297));
  INX1 g51682(.A (n_291), .Q (n_292));
  INX1 g51683(.A (n_290), .Q (n_289));
  INX1 g51684(.A (n_286), .Q (n_285));
  INX1 g51685(.A (n_284), .Q (n_283));
  INX1 g51686(.A (n_281), .Q (n_280));
  INX1 g51687(.A (n_279), .Q (n_278));
  INX1 g51688(.A (n_128), .Q (n_276));
  INX1 g51689(.A (n_275), .Q (n_274));
  INX1 g51690(.A (n_127), .Q (n_273));
  INX1 g51691(.A (n_272), .Q (n_271));
  AND2X1 g51693(.A (n_4534), .B (n_122), .Q (n_269));
  AND2X1 g51696(.A (n_5985), .B (n_121), .Q (n_268));
  AND2X1 g51702(.A (n_5730), .B (n_121), .Q (n_267));
  AND2X1 g51712(.A (n_4536), .B (n_121), .Q (n_266));
  AND2X1 g51719(.A (n_5749), .B (n_121), .Q (n_265));
  AND2X1 g51722(.A (n_5741), .B (n_121), .Q (n_264));
  AND2X1 g51726(.A (n_5748), .B (n_121), .Q (n_263));
  AND2X1 g51735(.A (n_5732), .B (n_121), .Q (n_262));
  AND2X1 g51737(.A (n_5736), .B (n_121), .Q (n_261));
  AND2X1 g51758(.A (n_5747), .B (n_122), .Q (n_260));
  AND2X1 g51771(.A (n_5738), .B (n_121), .Q (n_259));
  AND2X1 g51772(.A (n_5739), .B (n_121), .Q (n_258));
  AND2X1 g51778(.A (n_4534), .B (n_121), .Q (n_257));
  NO2X1 g51779(.A (alu_2nd_operand[1]), .B (n_6629), .Q (n_256));
  AND2X1 g51780(.A (n_5751), .B (n_122), .Q (n_255));
  AND2X1 g51793(.A (n_6731), .B (n_121), .Q (n_254));
  AND2X1 g51795(.A (n_5750), .B (n_122), .Q (n_253));
  AND2X1 g51798(.A (instruction[17]), .B (n_121), .Q (n_252));
  AND2X1 g51799(.A (instruction[15]), .B (n_121), .Q (n_251));
  AND2X1 g51800(.A (instruction[16]), .B (n_121), .Q (n_250));
  AND2X1 g51801(.A (instruction[18]), .B (n_121), .Q (n_249));
  AND2X1 g51802(.A (n_6723), .B (n_122), .Q (n_248));
  AND2X1 g51803(.A (instruction[21]), .B (n_122), .Q (n_247));
  AND2X1 g51804(.A (instruction[19]), .B (n_121), .Q (n_246));
  AND2X1 g51805(.A (instruction[23]), .B (n_121), .Q (n_245));
  AND2X1 g51806(.A (instruction[22]), .B (n_122), .Q (n_244));
  AND2X1 g51807(.A (instruction[24]), .B (n_122), .Q (n_243));
  AND2X1 g51808(.A (\instruction[5]_40139 ), .B (n_121), .Q (n_242));
  OR2X1 g51809(.A (n_6718), .B (n_123), .Q (n_241));
  OR2X1 g51810(.A (instruction[4]), .B (n_123), .Q (n_240));
  OR2X1 g51811(.A (instruction[0]), .B (n_123), .Q (n_239));
  AND2X1 g51812(.A (instruction[2]), .B (n_121), .Q (n_238));
  AND2X1 g51813(.A (instruction[3]), .B (n_121), .Q (n_237));
  NO2X1 g51814(.A (alu_2nd_operand[31]), .B (alu_sra_result[31]), .Q
       (n_236));
  NO2X1 g51815(.A (alu_2nd_operand[29]), .B (\rs1_data[29]_39336 ), .Q
       (n_235));
  AND2X1 g51816(.A (instruction[6]), .B (n_121), .Q (n_234));
  AND2X1 g51817(.A (n_6721), .B (n_121), .Q (n_233));
  AND2X1 g51818(.A (\instruction[7]_39562 ), .B (n_121), .Q (n_232));
  AND2X1 g51819(.A (n_6720), .B (n_122), .Q (n_231));
  AND2X1 g51820(.A (instruction[25]), .B (n_122), .Q (n_230));
  NO2X1 g51821(.A (alu_2nd_operand[20]), .B (n_4486), .Q (n_229));
  AND2X1 g51822(.A (\instruction[10]_39951 ), .B (n_121), .Q (n_228));
  AND2X1 g51823(.A (\instruction[11]_40800 ), .B (n_121), .Q (n_227));
  NO2X1 g51824(.A (n_178), .B (\rs1_data[0]_39306 ), .Q (n_226));
  AND2X1 g51825(.A (instruction[26]), .B (n_121), .Q (n_225));
  AND2X1 g51826(.A (\instruction[9]_39983 ), .B (n_121), .Q (n_224));
  AND2X1 g51827(.A (instruction[27]), .B (n_121), .Q (n_223));
  NO2X1 g51828(.A (alu_2nd_operand[21]), .B (n_4479), .Q (n_222));
  AND2X1 g51829(.A (\instruction[14]_40077 ), .B (n_122), .Q (n_221));
  AND2X1 g51830(.A (instruction[28]), .B (n_122), .Q (n_220));
  AND2X1 g51831(.A (n_6722), .B (n_122), .Q (n_219));
  AND2X1 g51832(.A (n_6719), .B (n_121), .Q (n_218));
  NO2X1 g51833(.A (alu_2nd_operand[22]), .B (n_4463), .Q (n_217));
  AND2X1 g51834(.A (\instruction[8]_40015 ), .B (n_122), .Q (n_216));
  NO2X1 g51835(.A (alu_2nd_operand[17]), .B (n_4482), .Q (n_215));
  AND2X1 g51836(.A (instruction[29]), .B (n_121), .Q (n_214));
  NO2X1 g51837(.A (alu_2nd_operand[23]), .B (\rs1_data[23]_39246 ), .Q
       (n_213));
  NA2I1X1 g51838(.B (n_4479), .AN (alu_2nd_operand[21]), .Q (n_341));
  OR2X1 g51839(.A (n_207), .B (n_4484), .Q (n_340));
  NA2X1 g51840(.A (n_210), .B (\rs1_data[14]_39466 ), .Q (n_339));
  NO2X1 g51842(.A (alu_2nd_operand[13]), .B (n_193), .Q (n_338));
  NO2X1 g51843(.A (alu_2nd_operand[12]), .B (n_192), .Q (n_336));
  NA2X1 g51844(.A (alu_2nd_operand[1]), .B (n_203), .Q (n_334));
  AND2X1 g51845(.A (n_178), .B (\rs1_data[0]_39306 ), .Q (n_333));
  NO2I1X1 g51846(.B (alu_2nd_operand[19]), .AN (n_4477), .Q (n_332));
  NA2I1X1 g51847(.B (\rs1_data[23]_39246 ), .AN (alu_2nd_operand[23]),
       .Q (n_331));
  NO2I1X1 g51848(.B (n_4478), .AN (alu_2nd_operand[18]), .Q (n_330));
  NO2X1 g51849(.A (n_4533), .B (\rs1_data[0]_39306 ), .Q (n_329));
  NO2X1 g51850(.A (n_177), .B (n_6757), .Q (n_328));
  OR2X1 g51851(.A (alu_2nd_operand[5]), .B (n_184), .Q (n_327));
  NO2X1 g51852(.A (alu_2nd_operand[6]), .B (n_187), .Q (n_326));
  NO2X1 g51853(.A (alu_2nd_operand[7]), .B (n_196), .Q (n_325));
  OR2X1 g51854(.A (alu_2nd_operand[15]), .B (n_188), .Q (n_324));
  NO2I1X1 g51855(.B (alu_2nd_operand[18]), .AN (n_4478), .Q (n_323));
  OR2X1 g51856(.A (alu_2nd_operand[31]), .B (n_198), .Q (n_322));
  OR2X1 g51857(.A (alu_2nd_operand[29]), .B (n_185), .Q (n_321));
  NA2I1X1 g51859(.B (n_4486), .AN (alu_2nd_operand[20]), .Q (n_320));
  NA2X1 g51860(.A (n_180), .B (n_4465), .Q (n_319));
  NO2I1X1 g51861(.B (alu_2nd_operand[17]), .AN (n_4482), .Q (n_318));
  NA2I1X1 g51862(.B (n_4463), .AN (alu_2nd_operand[22]), .Q (n_317));
  NO2I1X1 g51863(.B (n_4463), .AN (alu_2nd_operand[22]), .Q (n_315));
  NO2I1X1 g51864(.B (n_4479), .AN (alu_2nd_operand[21]), .Q (n_313));
  NA2X1 g51865(.A (alu_2nd_operand[25]), .B (n_199), .Q (n_311));
  NO2X1 g51866(.A (alu_2nd_operand[4]), .B (alu_2nd_operand[3]), .Q
       (n_310));
  NO2I1X1 g51867(.B (n_4482), .AN (alu_2nd_operand[17]), .Q (n_309));
  NA2X1 g51868(.A (alu_2nd_operand[11]), .B (n_202), .Q (n_307));
  NO2I1X1 g51869(.B (n_4477), .AN (alu_2nd_operand[19]), .Q (n_305));
  NA2X1 g51870(.A (alu_2nd_operand[27]), .B (n_194), .Q (n_304));
  NA2X1 g51871(.A (alu_2nd_operand[29]), .B (n_185), .Q (n_302));
  NA2X1 g51872(.A (alu_2nd_operand[31]), .B (n_198), .Q (n_300));
  NO2X1 g51873(.A (n_176), .B (n_6071), .Q (n_298));
  NA2X1 g51874(.A (alu_2nd_operand[9]), .B (n_200), .Q (n_296));
  NO2I1X1 g51875(.B (\rs1_data[23]_39246 ), .AN (alu_2nd_operand[23]),
       .Q (n_295));
  NO2X1 g51876(.A (n_180), .B (alu_2nd_operand[3]), .Q (n_294));
  NA2X1 g51877(.A (n_179), .B (n_6629), .Q (n_293));
  NA2X1 g51878(.A (n_179), .B (alu_2nd_operand[2]), .Q (n_291));
  NA2X1 g51879(.A (n_124), .B (alu_2nd_operand[3]), .Q (n_290));
  NO2X1 g51880(.A (alu_2nd_operand[1]), .B (alu_2nd_operand[2]), .Q
       (n_288));
  AND2X1 g51881(.A (n_201), .B (n_5605), .Q (n_287));
  NO2X1 g51882(.A (n_178), .B (n_198), .Q (n_286));
  NA2X1 g51883(.A (alu_2nd_operand[2]), .B (n_177), .Q (n_284));
  NO2X1 g51884(.A (alu_2nd_operand[4]), .B (n_177), .Q (n_282));
  AND2X1 g51885(.A (n_4533), .B (\rs1_data[0]_39306 ), .Q (n_281));
  NA2X1 g51886(.A (n_124), .B (n_177), .Q (n_279));
  AND2X1 g51887(.A (n_201), .B (n_6721), .Q (n_277));
  AND2X1 g51889(.A (n_179), .B (n_178), .Q (n_275));
  AND2X1 g51891(.A (alu_2nd_operand[1]), .B (n_178), .Q (n_272));
  NO2X1 g51892(.A (n_6601), .B (n_6600), .Q (n_270));
  INX1 g51895(.A (n_6067), .Q (n_212));
  INX1 g51903(.A (alu_2nd_operand[14]), .Q (n_210));
  INX1 g51907(.A (alu_2nd_operand[28]), .Q (n_209));
  INX1 g51908(.A (alu_2nd_operand[9]), .Q (n_208));
  INX1 g51909(.A (alu_2nd_operand[16]), .Q (n_207));
  INX1 g51910(.A (alu_2nd_operand[11]), .Q (n_206));
  INX1 g51911(.A (n_6726), .Q (n_205));
  INX1 g51913(.A (n_6629), .Q (n_203));
  INX1 g51914(.A (n_4474), .Q (n_202));
  INX1 g51916(.A (n_4487), .Q (n_200));
  INX1 g51917(.A (n_4481), .Q (n_199));
  INX1 g51918(.A (alu_sra_result[31]), .Q (n_198));
  INX1 g51920(.A (\rs1_data[14]_39466 ), .Q (n_197));
  INX1 g51921(.A (n_4460), .Q (n_196));
  INX1 g51922(.A (n_4480), .Q (n_195));
  INX1 g51923(.A (\rs1_data[27]_39286 ), .Q (n_194));
  INX1 g51924(.A (n_4476), .Q (n_193));
  INX1 g51925(.A (n_4475), .Q (n_192));
  INX1 g51927(.A (n_4464), .Q (n_190));
  INX1 g51929(.A (n_4483), .Q (n_189));
  INX1 g51930(.A (\rs1_data[15]_39476 ), .Q (n_188));
  INX1 g51931(.A (n_4466), .Q (n_187));
  INX1 g51932(.A (n_4485), .Q (n_186));
  INX1 g51933(.A (\rs1_data[29]_39336 ), .Q (n_185));
  INX1 g51934(.A (n_4461), .Q (n_184));
  INX1 g51935(.A (n_4465), .Q (n_183));
  INX1 g51936(.A (\rs1_data[26]_39276 ), .Q (n_182));
  INX1 g51937(.A (\rs1_data[28]_39296 ), .Q (n_181));
  INX1 g51939(.A (alu_2nd_operand[4]), .Q (n_180));
  INX1 g51940(.A (alu_2nd_operand[1]), .Q (n_179));
  INX1 g51941(.A (n_4533), .Q (n_178));
  INX1 g51943(.A (n_6453), .Q (n_176));
  INX1 g51955(.A (read_data[23]), .Q (n_174));
  INX1 g51970(.A (read_data[31]), .Q (n_173));
  DFRQX1 csr_mcause_interrupt_flag_reg(.C (rc_gclk_205603), .D (n_782),
       .Q (csr_mcause_interrupt_flag));
  DFRQX1 \csr_mcycle_reg[0] (.C (clock), .D (n_1155), .Q
       (csr_mcycle[0]));
  DFRQX1 \csr_mcycle_reg[10] (.C (clock), .D (n_1186), .Q
       (csr_mcycle[10]));
  DFRQX1 \csr_mcycle_reg[11] (.C (clock), .D (n_1190), .Q
       (csr_mcycle[11]));
  DFRQX1 \csr_mcycle_reg[12] (.C (clock), .D (n_1182), .Q
       (csr_mcycle[12]));
  DFRQX1 \csr_mcycle_reg[13] (.C (clock), .D (n_1185), .Q
       (csr_mcycle[13]));
  DFRQX1 \csr_mcycle_reg[14] (.C (clock), .D (n_1189), .Q
       (csr_mcycle[14]));
  DFRQX1 \csr_mcycle_reg[15] (.C (clock), .D (n_1194), .Q
       (csr_mcycle[15]));
  DFRQX1 \csr_mcycle_reg[16] (.C (clock), .D (n_1193), .Q
       (csr_mcycle[16]));
  DFRQX1 \csr_mcycle_reg[17] (.C (clock), .D (n_1199), .Q
       (csr_mcycle[17]));
  DFRQX1 \csr_mcycle_reg[18] (.C (clock), .D (n_1206), .Q
       (csr_mcycle[18]));
  DFRQX1 \csr_mcycle_reg[19] (.C (clock), .D (n_1219), .Q
       (csr_mcycle[19]));
  DFRQX1 \csr_mcycle_reg[1] (.C (clock), .D (n_1156), .Q
       (csr_mcycle[1]));
  DFRQX1 \csr_mcycle_reg[20] (.C (clock), .D (n_1198), .Q
       (csr_mcycle[20]));
  DFRQX1 \csr_mcycle_reg[21] (.C (clock), .D (n_1205), .Q
       (csr_mcycle[21]));
  DFRQX1 \csr_mcycle_reg[22] (.C (clock), .D (n_1221), .Q
       (csr_mcycle[22]));
  DFRQX1 \csr_mcycle_reg[23] (.C (clock), .D (n_1228), .Q
       (csr_mcycle[23]));
  DFRQX1 \csr_mcycle_reg[24] (.C (clock), .D (n_1197), .Q
       (csr_mcycle[24]));
  DFRQX1 \csr_mcycle_reg[25] (.C (clock), .D (n_1204), .Q
       (csr_mcycle[25]));
  DFRQX1 \csr_mcycle_reg[26] (.C (clock), .D (n_1220), .Q
       (csr_mcycle[26]));
  DFRQX1 \csr_mcycle_reg[27] (.C (clock), .D (n_1227), .Q
       (csr_mcycle[27]));
  DFRQX1 \csr_mcycle_reg[28] (.C (clock), .D (n_1207), .Q
       (csr_mcycle[28]));
  DFRQX1 \csr_mcycle_reg[29] (.C (clock), .D (n_1222), .Q
       (csr_mcycle[29]));
  DFRQX1 \csr_mcycle_reg[2] (.C (clock), .D (n_1161), .Q
       (csr_mcycle[2]));
  DFRQX1 \csr_mcycle_reg[30] (.C (clock), .D (n_1226), .Q
       (csr_mcycle[30]));
  DFRQX1 \csr_mcycle_reg[31] (.C (clock), .D (n_1231), .Q
       (csr_mcycle[31]));
  DFRQX1 \csr_mcycle_reg[35] (.C (clock), .D (n_1249), .Q
       (csr_mcycle[35]));
  DFRQX1 \csr_mcycle_reg[39] (.C (clock), .D (n_1257), .Q
       (csr_mcycle[39]));
  DFRQX1 \csr_mcycle_reg[3] (.C (clock), .D (n_1166), .Q
       (csr_mcycle[3]));
  DFRQX1 \csr_mcycle_reg[43] (.C (clock), .D (n_1268), .Q
       (csr_mcycle[43]));
  DFRQX1 \csr_mcycle_reg[47] (.C (clock), .D (n_1276), .Q
       (csr_mcycle[47]));
  DFRQX1 \csr_mcycle_reg[4] (.C (clock), .D (n_1167), .Q
       (csr_mcycle[4]));
  DFRQX1 \csr_mcycle_reg[51] (.C (clock), .D (n_1275), .Q
       (csr_mcycle[51]));
  DFRQX1 \csr_mcycle_reg[55] (.C (clock), .D (n_1285), .Q
       (csr_mcycle[55]));
  DFRQX2 \csr_mcycle_reg[56] (.C (clock), .D (n_1273), .Q
       (csr_mcycle[56]));
  DFRQX2 \csr_mcycle_reg[58] (.C (clock), .D (n_1286), .Q
       (csr_mcycle[58]));
  DFRQX1 \csr_mcycle_reg[59] (.C (clock), .D (n_1291), .Q
       (csr_mcycle[59]));
  DFRQX1 \csr_mcycle_reg[5] (.C (clock), .D (n_1173), .Q
       (csr_mcycle[5]));
  DFRQX1 \csr_mcycle_reg[60] (.C (clock), .D (n_1279), .Q
       (csr_mcycle[60]));
  DFRQX1 \csr_mcycle_reg[62] (.C (clock), .D (n_1292), .Q
       (csr_mcycle[62]));
  DFRQX1 \csr_mcycle_reg[63] (.C (clock), .D (n_1293), .Q
       (csr_mcycle[63]));
  DFRQX1 \csr_mcycle_reg[6] (.C (clock), .D (n_1175), .Q
       (csr_mcycle[6]));
  DFRQX1 \csr_mcycle_reg[7] (.C (clock), .D (n_1177), .Q
       (csr_mcycle[7]));
  DFRQX1 \csr_mcycle_reg[8] (.C (clock), .D (n_1178), .Q
       (csr_mcycle[8]));
  DFRQX1 \csr_mcycle_reg[9] (.C (clock), .D (n_1181), .Q
       (csr_mcycle[9]));
  DFRQX1 \csr_mepc_reg[10] (.C (rc_gclk_205556), .D (n_781), .Q
       (n_5557));
  DFRQX1 \csr_mepc_reg[11] (.C (rc_gclk_205556), .D (n_772), .Q
       (n_5556));
  DFRQX1 \csr_mepc_reg[12] (.C (rc_gclk_205556), .D (n_760), .Q
       (n_5555));
  DFRQX1 \csr_mepc_reg[13] (.C (rc_gclk_205556), .D (n_759), .Q
       (n_5553));
  DFRQX1 \csr_mepc_reg[14] (.C (rc_gclk_205556), .D (n_778), .Q
       (n_5552));
  DFRQX1 \csr_mepc_reg[15] (.C (rc_gclk_205556), .D (n_777), .Q
       (n_5551));
  DFRQX1 \csr_mepc_reg[16] (.C (rc_gclk_205556), .D (n_771), .Q
       (n_5550));
  DFRQX1 \csr_mepc_reg[17] (.C (rc_gclk_205556), .D (n_770), .Q
       (n_5549));
  DFRQX1 \csr_mepc_reg[18] (.C (rc_gclk_205556), .D (n_769), .Q
       (n_5548));
  DFRQX1 \csr_mepc_reg[19] (.C (rc_gclk_205556), .D (n_758), .Q
       (n_5547));
  DFRQX1 \csr_mepc_reg[20] (.C (rc_gclk_205556), .D (n_757), .Q
       (n_5546));
  DFRQX1 \csr_mepc_reg[21] (.C (rc_gclk_205556), .D (n_756), .Q
       (n_5545));
  DFRQX1 \csr_mepc_reg[22] (.C (rc_gclk_205556), .D (n_768), .Q
       (n_5544));
  DFRQX1 \csr_mepc_reg[23] (.C (rc_gclk_205556), .D (n_767), .Q
       (n_5572));
  DFRQX1 \csr_mepc_reg[24] (.C (rc_gclk_205556), .D (n_755), .Q
       (n_5571));
  DFRQX1 \csr_mepc_reg[25] (.C (rc_gclk_205556), .D (n_754), .Q
       (n_5570));
  DFRQX1 \csr_mepc_reg[26] (.C (rc_gclk_205556), .D (n_776), .Q
       (n_5569));
  DFRQX1 \csr_mepc_reg[27] (.C (rc_gclk_205556), .D (n_766), .Q
       (n_5568));
  DFRQX1 \csr_mepc_reg[28] (.C (rc_gclk_205556), .D (n_775), .Q
       (n_5567));
  DFRQX1 \csr_mepc_reg[29] (.C (rc_gclk_205556), .D (n_774), .Q
       (n_5565));
  DFRQX1 \csr_mepc_reg[2] (.C (rc_gclk_205556), .D (n_765), .Q
       (n_5566));
  DFRQX1 \csr_mepc_reg[30] (.C (rc_gclk_205556), .D (n_773), .Q
       (n_5554));
  DFRQX1 \csr_mepc_reg[31] (.C (rc_gclk_205556), .D (n_780), .Q
       (n_5543));
  DFRQX1 \csr_mepc_reg[3] (.C (rc_gclk_205556), .D (n_764), .Q
       (n_5564));
  DFRQX1 \csr_mepc_reg[4] (.C (rc_gclk_205556), .D (n_779), .Q
       (n_5563));
  DFRQX1 \csr_mepc_reg[5] (.C (rc_gclk_205556), .D (n_763), .Q
       (n_5562));
  DFRQX1 \csr_mepc_reg[6] (.C (rc_gclk_205556), .D (n_753), .Q
       (n_5561));
  DFRQX1 \csr_mepc_reg[7] (.C (rc_gclk_205556), .D (n_752), .Q
       (n_5560));
  DFRQX1 \csr_mepc_reg[8] (.C (rc_gclk_205556), .D (n_761), .Q
       (n_5559));
  DFRQX1 \csr_mepc_reg[9] (.C (rc_gclk_205556), .D (n_762), .Q
       (n_5558));
  DFRQX1 csr_mie_meie_reg(.C (rc_gclk_205601), .D (n_104), .Q (n_6322));
  DFRQX1 \csr_mie_mfie_reg[0] (.C (rc_gclk_205601), .D (n_101), .Q
       (n_6326));
  DFRQX1 \csr_mie_mfie_reg[10] (.C (rc_gclk_205601), .D (n_81), .Q
       (n_6338));
  DFRQX1 \csr_mie_mfie_reg[11] (.C (rc_gclk_205601), .D (n_95), .Q
       (n_6339));
  DFRQX1 \csr_mie_mfie_reg[12] (.C (rc_gclk_205601), .D (n_82), .Q
       (n_6340));
  DFRQX1 \csr_mie_mfie_reg[13] (.C (rc_gclk_205601), .D (n_94), .Q
       (n_6342));
  DFRQX1 \csr_mie_mfie_reg[14] (.C (rc_gclk_205601), .D (n_83), .Q
       (n_6343));
  DFRQX1 \csr_mie_mfie_reg[15] (.C (rc_gclk_205601), .D (n_84), .Q
       (n_6344));
  DFRQX1 \csr_mie_mfie_reg[1] (.C (rc_gclk_205601), .D (n_100), .Q
       (n_6327));
  DFRQX1 \csr_mie_mfie_reg[2] (.C (rc_gclk_205601), .D (n_99), .Q
       (n_6328));
  DFRQX1 \csr_mie_mfie_reg[3] (.C (rc_gclk_205601), .D (n_98), .Q
       (n_6330));
  DFRQX1 \csr_mie_mfie_reg[4] (.C (rc_gclk_205601), .D (n_89), .Q
       (n_6331));
  DFRQX1 \csr_mie_mfie_reg[5] (.C (rc_gclk_205601), .D (n_97), .Q
       (n_6332));
  DFRQX1 \csr_mie_mfie_reg[6] (.C (rc_gclk_205601), .D (n_79), .Q
       (n_6333));
  DFRQX1 \csr_mie_mfie_reg[7] (.C (rc_gclk_205601), .D (n_88), .Q
       (n_6334));
  DFRQX1 \csr_mie_mfie_reg[8] (.C (rc_gclk_205601), .D (n_96), .Q
       (n_6336));
  DFRQX1 \csr_mie_mfie_reg[9] (.C (rc_gclk_205601), .D (n_80), .Q
       (n_6337));
  DFRQX1 csr_mie_msie_reg(.C (rc_gclk_205601), .D (n_86), .Q (n_6325));
  DFRQX1 csr_mie_mtie_reg(.C (rc_gclk_205601), .D (n_105), .Q (n_6324));
  DFRQX1 \csr_minstret_reg[0] (.C (rc_gclk), .D (n_1157), .Q
       (csr_minstret[0]));
  DFRQX1 \csr_minstret_reg[10] (.C (rc_gclk), .D (n_1187), .Q
       (csr_minstret[10]));
  DFRQX1 \csr_minstret_reg[11] (.C (rc_gclk), .D (n_1191), .Q
       (csr_minstret[11]));
  DFRQX1 \csr_minstret_reg[12] (.C (rc_gclk), .D (n_1184), .Q
       (csr_minstret[12]));
  DFRQX1 \csr_minstret_reg[13] (.C (rc_gclk), .D (n_1188), .Q
       (csr_minstret[13]));
  DFRQX1 \csr_minstret_reg[14] (.C (rc_gclk), .D (n_1192), .Q
       (csr_minstret[14]));
  DFRQX1 \csr_minstret_reg[15] (.C (rc_gclk), .D (n_1196), .Q
       (csr_minstret[15]));
  DFRQX2 \csr_minstret_reg[18] (.C (rc_gclk), .D (n_1216), .Q
       (csr_minstret[18]));
  DFRQX1 \csr_minstret_reg[19] (.C (rc_gclk), .D (n_1224), .Q
       (csr_minstret[19]));
  DFRQX1 \csr_minstret_reg[1] (.C (rc_gclk), .D (n_1160), .Q
       (csr_minstret[1]));
  DFRQX1 \csr_minstret_reg[21] (.C (rc_gclk), .D (n_1169), .Q
       (csr_minstret[21]));
  DFRQX1 \csr_minstret_reg[22] (.C (rc_gclk), .D (n_1203), .Q
       (csr_minstret[22]));
  DFRQX1 \csr_minstret_reg[23] (.C (rc_gclk), .D (n_1218), .Q
       (csr_minstret[23]));
  DFRQX1 \csr_minstret_reg[24] (.C (rc_gclk), .D (n_1200), .Q
       (csr_minstret[24]));
  DFRQX1 \csr_minstret_reg[25] (.C (rc_gclk), .D (n_1208), .Q
       (csr_minstret[25]));
  DFRQX1 \csr_minstret_reg[26] (.C (rc_gclk), .D (n_1223), .Q
       (csr_minstret[26]));
  DFRQX1 \csr_minstret_reg[27] (.C (rc_gclk), .D (n_1229), .Q
       (csr_minstret[27]));
  DFRQX1 \csr_minstret_reg[28] (.C (rc_gclk), .D (n_1217), .Q
       (csr_minstret[28]));
  DFRQX1 \csr_minstret_reg[29] (.C (rc_gclk), .D (n_1225), .Q
       (csr_minstret[29]));
  DFRQX1 \csr_minstret_reg[2] (.C (rc_gclk), .D (n_1165), .Q
       (csr_minstret[2]));
  DFRQX2 \csr_minstret_reg[30] (.C (rc_gclk), .D (n_1230), .Q
       (csr_minstret[30]));
  DFRQX1 \csr_minstret_reg[31] (.C (rc_gclk), .D (n_1232), .Q
       (csr_minstret[31]));
  DFRQX2 \csr_minstret_reg[33] (.C (rc_gclk), .D (n_1238), .Q
       (csr_minstret[33]));
  DFRQX2 \csr_minstret_reg[34] (.C (rc_gclk), .D (n_1242), .Q
       (csr_minstret[34]));
  DFRQX1 \csr_minstret_reg[35] (.C (rc_gclk), .D (n_1252), .Q
       (csr_minstret[35]));
  DFRQX2 \csr_minstret_reg[36] (.C (rc_gclk), .D (n_1237), .Q
       (csr_minstret[36]));
  DFRQX2 \csr_minstret_reg[37] (.C (rc_gclk), .D (n_1243), .Q
       (csr_minstret[37]));
  DFRQX1 \csr_minstret_reg[39] (.C (rc_gclk), .D (n_1264), .Q
       (csr_minstret[39]));
  DFRQX1 \csr_minstret_reg[3] (.C (rc_gclk), .D (n_1170), .Q
       (csr_minstret[3]));
  DFRQX1 \csr_minstret_reg[43] (.C (rc_gclk), .D (n_1272), .Q
       (csr_minstret[43]));
  DFRQX2 \csr_minstret_reg[44] (.C (rc_gclk), .D (n_1253), .Q
       (csr_minstret[44]));
  DFRQX2 \csr_minstret_reg[45] (.C (rc_gclk), .D (n_1262), .Q
       (csr_minstret[45]));
  DFRQX2 \csr_minstret_reg[46] (.C (rc_gclk), .D (n_1271), .Q
       (csr_minstret[46]));
  DFRQX1 \csr_minstret_reg[47] (.C (rc_gclk), .D (n_1282), .Q
       (csr_minstret[47]));
  DFRQX2 \csr_minstret_reg[48] (.C (rc_gclk), .D (n_1251), .Q
       (csr_minstret[48]));
  DFRQX2 \csr_minstret_reg[49] (.C (rc_gclk), .D (n_1261), .Q
       (csr_minstret[49]));
  DFRQX1 \csr_minstret_reg[4] (.C (rc_gclk), .D (n_1172), .Q
       (csr_minstret[4]));
  DFRQX1 \csr_minstret_reg[51] (.C (rc_gclk), .D (n_1281), .Q
       (csr_minstret[51]));
  DFRQX2 \csr_minstret_reg[52] (.C (rc_gclk), .D (n_1260), .Q
       (csr_minstret[52]));
  DFRQX2 \csr_minstret_reg[54] (.C (rc_gclk), .D (n_1280), .Q
       (csr_minstret[54]));
  DFRQX1 \csr_minstret_reg[55] (.C (rc_gclk), .D (n_1287), .Q
       (csr_minstret[55]));
  DFRQX2 \csr_minstret_reg[56] (.C (rc_gclk), .D (n_1277), .Q
       (csr_minstret[56]));
  DFRQX2 \csr_minstret_reg[57] (.C (rc_gclk), .D (n_1283), .Q
       (csr_minstret[57]));
  DFRQX2 \csr_minstret_reg[58] (.C (rc_gclk), .D (n_1288), .Q
       (csr_minstret[58]));
  DFRQX1 \csr_minstret_reg[59] (.C (rc_gclk), .D (n_1294), .Q
       (csr_minstret[59]));
  DFRQX1 \csr_minstret_reg[5] (.C (rc_gclk), .D (n_1174), .Q
       (csr_minstret[5]));
  DFRQX1 \csr_minstret_reg[60] (.C (rc_gclk), .D (n_1284), .Q
       (csr_minstret[60]));
  DFRQX2 \csr_minstret_reg[61] (.C (rc_gclk), .D (n_1290), .Q
       (csr_minstret[61]));
  DFRQX1 \csr_minstret_reg[62] (.C (rc_gclk), .D (n_1256), .Q
       (csr_minstret[62]));
  DFRQX1 \csr_minstret_reg[63] (.C (rc_gclk), .D (n_1295), .Q
       (csr_minstret[63]));
  DFRQX2 \csr_minstret_reg[6] (.C (rc_gclk), .D (n_1176), .Q
       (csr_minstret[6]));
  DFRQX1 \csr_minstret_reg[7] (.C (rc_gclk), .D (n_1179), .Q
       (csr_minstret[7]));
  DFRQX1 \csr_minstret_reg[8] (.C (rc_gclk), .D (n_1180), .Q
       (csr_minstret[8]));
  DFRQX1 \csr_minstret_reg[9] (.C (rc_gclk), .D (n_1183), .Q
       (csr_minstret[9]));
  DFRQX1 \csr_mtvec_reg[0] (.C (rc_gclk_205598), .D (n_269), .Q
       (n_6345));
  DFRQX1 \csr_mtvec_reg[10] (.C (rc_gclk_205598), .D (n_91), .Q
       (csr_mtvec[10]));
  DFRQX1 \csr_mtvec_reg[11] (.C (rc_gclk_205598), .D (n_104), .Q
       (csr_mtvec[11]));
  DFRQX1 \csr_mtvec_reg[12] (.C (rc_gclk_205598), .D (n_260), .Q
       (csr_mtvec[12]));
  DFRQX1 \csr_mtvec_reg[13] (.C (rc_gclk_205598), .D (n_103), .Q
       (csr_mtvec[13]));
  DFRQX1 \csr_mtvec_reg[14] (.C (rc_gclk_205598), .D (n_90), .Q
       (csr_mtvec[14]));
  DFRQX1 \csr_mtvec_reg[15] (.C (rc_gclk_205598), .D (n_102), .Q
       (csr_mtvec[15]));
  DFRQX1 \csr_mtvec_reg[16] (.C (rc_gclk_205598), .D (n_101), .Q
       (csr_mtvec[16]));
  DFRQX1 \csr_mtvec_reg[17] (.C (rc_gclk_205598), .D (n_100), .Q
       (csr_mtvec[17]));
  DFRQX1 \csr_mtvec_reg[18] (.C (rc_gclk_205598), .D (n_99), .Q
       (csr_mtvec[18]));
  DFRQX1 \csr_mtvec_reg[19] (.C (rc_gclk_205598), .D (n_98), .Q
       (csr_mtvec[19]));
  DFRQX1 \csr_mtvec_reg[20] (.C (rc_gclk_205598), .D (n_89), .Q
       (csr_mtvec[20]));
  DFRQX1 \csr_mtvec_reg[21] (.C (rc_gclk_205598), .D (n_97), .Q
       (csr_mtvec[21]));
  DFRQX1 \csr_mtvec_reg[22] (.C (rc_gclk_205598), .D (n_79), .Q
       (csr_mtvec[22]));
  DFRQX1 \csr_mtvec_reg[23] (.C (rc_gclk_205598), .D (n_88), .Q
       (csr_mtvec[23]));
  DFRQX1 \csr_mtvec_reg[24] (.C (rc_gclk_205598), .D (n_96), .Q
       (csr_mtvec[24]));
  DFRQX1 \csr_mtvec_reg[25] (.C (rc_gclk_205598), .D (n_80), .Q
       (csr_mtvec[25]));
  DFRQX1 \csr_mtvec_reg[26] (.C (rc_gclk_205598), .D (n_81), .Q
       (csr_mtvec[26]));
  DFRQX1 \csr_mtvec_reg[27] (.C (rc_gclk_205598), .D (n_95), .Q
       (csr_mtvec[27]));
  DFRQX1 \csr_mtvec_reg[28] (.C (rc_gclk_205598), .D (n_82), .Q
       (csr_mtvec[28]));
  DFRQX1 \csr_mtvec_reg[29] (.C (rc_gclk_205598), .D (n_94), .Q
       (csr_mtvec[29]));
  DFRQX1 \csr_mtvec_reg[2] (.C (rc_gclk_205598), .D (n_87), .Q
       (csr_mtvec[2]));
  DFRQX1 \csr_mtvec_reg[30] (.C (rc_gclk_205598), .D (n_83), .Q
       (csr_mtvec[30]));
  DFRQX1 \csr_mtvec_reg[31] (.C (rc_gclk_205598), .D (n_84), .Q
       (csr_mtvec[31]));
  DFRQX1 \csr_mtvec_reg[3] (.C (rc_gclk_205598), .D (n_86), .Q
       (csr_mtvec[3]));
  DFRQX1 \csr_mtvec_reg[4] (.C (rc_gclk_205598), .D (n_85), .Q
       (csr_mtvec[4]));
  DFRQX1 \csr_mtvec_reg[5] (.C (rc_gclk_205598), .D (n_93), .Q
       (csr_mtvec[5]));
  DFRQX1 \csr_mtvec_reg[6] (.C (rc_gclk_205598), .D (n_92), .Q
       (csr_mtvec[6]));
  DFRQX1 \csr_mtvec_reg[7] (.C (rc_gclk_205598), .D (n_105), .Q
       (csr_mtvec[7]));
  DFRQX1 \csr_mtvec_reg[8] (.C (rc_gclk_205598), .D (n_255), .Q
       (csr_mtvec[8]));
  DFRQX1 \csr_mtvec_reg[9] (.C (rc_gclk_205598), .D (n_253), .Q
       (csr_mtvec[9]));
  DFRQX1 \current_state_reg[0] (.C (rc_gclk_205606), .D (n_123), .Q
       (current_state[0]));
  DFRQX1 \current_state_reg[1] (.C (rc_gclk_205606), .D (n_751), .Q
       (current_state[1]));
  DFRQX1 \current_state_reg[2] (.C (rc_gclk_205606), .D (n_564), .Q
       (current_state[2]));
  DFRQX1 \current_state_reg[3] (.C (rc_gclk_205606), .D (n_750), .Q
       (current_state[3]));
  DFRQX1 \integer_file_reg[10][0] (.C (rc_gclk_205535), .D (n_26), .Q
       (n_4757));
  DFRQX1 \integer_file_reg[10][10] (.C (rc_gclk_205535), .D (n_78), .Q
       (n_5098));
  DFRQX1 \integer_file_reg[10][11] (.C (rc_gclk_205535), .D (n_77), .Q
       (n_5129));
  DFRQX1 \integer_file_reg[10][12] (.C (rc_gclk_205535), .D (n_38), .Q
       (n_5160));
  DFRQX1 \integer_file_reg[10][13] (.C (rc_gclk_205535), .D (n_54), .Q
       (n_5222));
  DFRQX1 \integer_file_reg[10][14] (.C (rc_gclk_205535), .D (n_37), .Q
       (n_5253));
  DFRQX1 \integer_file_reg[10][15] (.C (rc_gclk_205535), .D (n_53), .Q
       (n_5284));
  DFRQX1 \integer_file_reg[10][16] (.C (rc_gclk_205535), .D (n_76), .Q
       (n_5315));
  DFRQX1 \integer_file_reg[10][17] (.C (rc_gclk_205535), .D (n_75), .Q
       (n_5346));
  DFRQX1 \integer_file_reg[10][18] (.C (rc_gclk_205535), .D (n_52), .Q
       (n_5377));
  DFRQX1 \integer_file_reg[10][19] (.C (rc_gclk_205535), .D (n_51), .Q
       (n_5408));
  DFRQX1 \integer_file_reg[10][1] (.C (rc_gclk_205535), .D (n_18), .Q
       (n_4788));
  DFRQX1 \integer_file_reg[10][20] (.C (rc_gclk_205535), .D (n_74), .Q
       (n_5439));
  DFRQX1 \integer_file_reg[10][21] (.C (rc_gclk_205535), .D (n_73), .Q
       (n_5470));
  DFRQX1 \integer_file_reg[10][22] (.C (rc_gclk_205535), .D (n_72), .Q
       (n_5501));
  DFRQX1 \integer_file_reg[10][23] (.C (rc_gclk_205535), .D (n_71), .Q
       (n_4571));
  DFRQX1 \integer_file_reg[10][24] (.C (rc_gclk_205535), .D (n_70), .Q
       (n_4602));
  DFRQX1 \integer_file_reg[10][25] (.C (rc_gclk_205535), .D (n_36), .Q
       (n_4633));
  DFRQX1 \integer_file_reg[10][26] (.C (rc_gclk_205535), .D (n_35), .Q
       (n_4664));
  DFRQX1 \integer_file_reg[10][27] (.C (rc_gclk_205535), .D (n_69), .Q
       (n_4695));
  DFRQX1 \integer_file_reg[10][28] (.C (rc_gclk_205535), .D (n_50), .Q
       (n_4726));
  DFRQX1 \integer_file_reg[10][29] (.C (rc_gclk_205535), .D (n_49), .Q
       (n_4850));
  DFRQX1 \integer_file_reg[10][2] (.C (rc_gclk_205535), .D (n_17), .Q
       (n_4819));
  DFRQX1 \integer_file_reg[10][30] (.C (rc_gclk_205535), .D (n_48), .Q
       (n_5191));
  DFRQX1 \integer_file_reg[10][31] (.C (rc_gclk_205535), .D (n_68), .Q
       (n_5532));
  DFRQX1 \integer_file_reg[10][3] (.C (rc_gclk_205535), .D (n_25), .Q
       (n_4881));
  DFRQX1 \integer_file_reg[10][4] (.C (rc_gclk_205535), .D (n_24), .Q
       (n_4912));
  DFRQX1 \integer_file_reg[10][5] (.C (rc_gclk_205535), .D (n_34), .Q
       (n_4943));
  DFRQX1 \integer_file_reg[10][6] (.C (rc_gclk_205535), .D (n_23), .Q
       (n_4974));
  DFRQX1 \integer_file_reg[10][7] (.C (rc_gclk_205535), .D (n_33), .Q
       (n_5005));
  DFRQX1 \integer_file_reg[10][8] (.C (rc_gclk_205535), .D (n_67), .Q
       (n_5036));
  DFRQX1 \integer_file_reg[10][9] (.C (rc_gclk_205535), .D (n_47), .Q
       (n_5067));
  DFRQX1 \integer_file_reg[11][0] (.C (rc_gclk_205559), .D (n_26), .Q
       (n_4756));
  DFRQX1 \integer_file_reg[11][10] (.C (rc_gclk_205559), .D (n_78), .Q
       (n_5097));
  DFRQX1 \integer_file_reg[11][11] (.C (rc_gclk_205559), .D (n_66), .Q
       (n_5128));
  DFRQX1 \integer_file_reg[11][12] (.C (rc_gclk_205559), .D (n_38), .Q
       (n_5159));
  DFRQX1 \integer_file_reg[11][13] (.C (rc_gclk_205559), .D (n_54), .Q
       (n_5221));
  DFRQX1 \integer_file_reg[11][14] (.C (rc_gclk_205559), .D (n_32), .Q
       (n_5252));
  DFRQX1 \integer_file_reg[11][15] (.C (rc_gclk_205559), .D (n_46), .Q
       (n_5283));
  DFRQX1 \integer_file_reg[11][16] (.C (rc_gclk_205559), .D (n_65), .Q
       (n_5314));
  DFRQX1 \integer_file_reg[11][17] (.C (rc_gclk_205559), .D (n_75), .Q
       (n_5345));
  DFRQX1 \integer_file_reg[11][18] (.C (rc_gclk_205559), .D (n_52), .Q
       (n_5376));
  DFRQX1 \integer_file_reg[11][19] (.C (rc_gclk_205559), .D (n_51), .Q
       (n_5407));
  DFRQX1 \integer_file_reg[11][1] (.C (rc_gclk_205559), .D (n_18), .Q
       (n_4787));
  DFRQX1 \integer_file_reg[11][20] (.C (rc_gclk_205559), .D (n_74), .Q
       (n_5438));
  DFRQX1 \integer_file_reg[11][21] (.C (rc_gclk_205559), .D (n_73), .Q
       (n_5469));
  DFRQX1 \integer_file_reg[11][22] (.C (rc_gclk_205559), .D (n_72), .Q
       (n_5500));
  DFRQX1 \integer_file_reg[11][23] (.C (rc_gclk_205559), .D (n_71), .Q
       (n_4570));
  DFRQX1 \integer_file_reg[11][24] (.C (rc_gclk_205559), .D (n_64), .Q
       (n_4601));
  DFRQX1 \integer_file_reg[11][25] (.C (rc_gclk_205559), .D (n_36), .Q
       (n_4632));
  DFRQX1 \integer_file_reg[11][26] (.C (rc_gclk_205559), .D (n_31), .Q
       (n_4663));
  DFRQX1 \integer_file_reg[11][27] (.C (rc_gclk_205559), .D (n_69), .Q
       (n_4694));
  DFRQX1 \integer_file_reg[11][28] (.C (rc_gclk_205559), .D (n_50), .Q
       (n_4725));
  DFRQX1 \integer_file_reg[11][29] (.C (rc_gclk_205559), .D (n_49), .Q
       (n_4849));
  DFRQX1 \integer_file_reg[11][2] (.C (rc_gclk_205559), .D (n_16), .Q
       (n_4818));
  DFRQX1 \integer_file_reg[11][30] (.C (rc_gclk_205559), .D (n_45), .Q
       (n_5190));
  DFRQX1 \integer_file_reg[11][31] (.C (rc_gclk_205559), .D (n_63), .Q
       (n_5531));
  DFRQX1 \integer_file_reg[11][3] (.C (rc_gclk_205559), .D (n_25), .Q
       (n_4880));
  DFRQX1 \integer_file_reg[11][4] (.C (rc_gclk_205559), .D (n_22), .Q
       (n_4911));
  DFRQX1 \integer_file_reg[11][5] (.C (rc_gclk_205559), .D (n_30), .Q
       (n_4942));
  DFRQX1 \integer_file_reg[11][6] (.C (rc_gclk_205559), .D (n_23), .Q
       (n_4973));
  DFRQX1 \integer_file_reg[11][7] (.C (rc_gclk_205559), .D (n_29), .Q
       (n_5004));
  DFRQX1 \integer_file_reg[11][8] (.C (rc_gclk_205559), .D (n_67), .Q
       (n_5035));
  DFRQX1 \integer_file_reg[11][9] (.C (rc_gclk_205559), .D (n_47), .Q
       (n_5066));
  DFRQX1 \integer_file_reg[12][0] (.C (rc_gclk_205568), .D (n_21), .Q
       (n_4755));
  DFRQX1 \integer_file_reg[12][10] (.C (rc_gclk_205568), .D (n_62), .Q
       (n_5096));
  DFRQX1 \integer_file_reg[12][11] (.C (rc_gclk_205568), .D (n_66), .Q
       (n_5127));
  DFRQX1 \integer_file_reg[12][12] (.C (rc_gclk_205568), .D (n_28), .Q
       (n_5158));
  DFRQX1 \integer_file_reg[12][13] (.C (rc_gclk_205568), .D (n_44), .Q
       (n_5220));
  DFRQX1 \integer_file_reg[12][14] (.C (rc_gclk_205568), .D (n_32), .Q
       (n_5251));
  DFRQX1 \integer_file_reg[12][15] (.C (rc_gclk_205568), .D (n_53), .Q
       (n_5282));
  DFRQX1 \integer_file_reg[12][16] (.C (rc_gclk_205568), .D (n_76), .Q
       (n_5313));
  DFRQX1 \integer_file_reg[12][17] (.C (rc_gclk_205568), .D (n_61), .Q
       (n_5344));
  DFRQX1 \integer_file_reg[12][18] (.C (rc_gclk_205568), .D (n_43), .Q
       (n_5375));
  DFRQX1 \integer_file_reg[12][19] (.C (rc_gclk_205568), .D (n_51), .Q
       (n_5406));
  DFRQX1 \integer_file_reg[12][1] (.C (rc_gclk_205568), .D (n_15), .Q
       (n_4786));
  DFRQX1 \integer_file_reg[12][20] (.C (rc_gclk_205568), .D (n_60), .Q
       (n_5437));
  DFRQX1 \integer_file_reg[12][21] (.C (rc_gclk_205568), .D (n_59), .Q
       (n_5468));
  DFRQX1 \integer_file_reg[12][22] (.C (rc_gclk_205568), .D (n_72), .Q
       (n_5499));
  DFRQX1 \integer_file_reg[12][23] (.C (rc_gclk_205568), .D (n_71), .Q
       (n_4569));
  DFRQX1 \integer_file_reg[12][24] (.C (rc_gclk_205568), .D (n_70), .Q
       (n_4600));
  DFRQX1 \integer_file_reg[12][25] (.C (rc_gclk_205568), .D (n_36), .Q
       (n_4631));
  DFRQX1 \integer_file_reg[12][26] (.C (rc_gclk_205568), .D (n_31), .Q
       (n_4662));
  DFRQX1 \integer_file_reg[12][27] (.C (rc_gclk_205568), .D (n_58), .Q
       (n_4693));
  DFRQX1 \integer_file_reg[12][28] (.C (rc_gclk_205568), .D (n_50), .Q
       (n_4724));
  DFRQX1 \integer_file_reg[12][29] (.C (rc_gclk_205568), .D (n_42), .Q
       (n_4848));
  DFRQX1 \integer_file_reg[12][2] (.C (rc_gclk_205568), .D (n_16), .Q
       (n_4817));
  DFRQX1 \integer_file_reg[12][30] (.C (rc_gclk_205568), .D (n_45), .Q
       (n_5189));
  DFRQX1 \integer_file_reg[12][31] (.C (rc_gclk_205568), .D (n_68), .Q
       (n_5530));
  DFRQX1 \integer_file_reg[12][3] (.C (rc_gclk_205568), .D (n_25), .Q
       (n_4879));
  DFRQX1 \integer_file_reg[12][4] (.C (rc_gclk_205568), .D (n_22), .Q
       (n_4910));
  DFRQX1 \integer_file_reg[12][5] (.C (rc_gclk_205568), .D (n_34), .Q
       (n_4941));
  DFRQX1 \integer_file_reg[12][6] (.C (rc_gclk_205568), .D (n_23), .Q
       (n_4972));
  DFRQX1 \integer_file_reg[12][7] (.C (rc_gclk_205568), .D (n_29), .Q
       (n_5003));
  DFRQX1 \integer_file_reg[12][8] (.C (rc_gclk_205568), .D (n_67), .Q
       (n_5034));
  DFRQX1 \integer_file_reg[12][9] (.C (rc_gclk_205568), .D (n_47), .Q
       (n_5065));
  DFRQX1 \integer_file_reg[13][0] (.C (rc_gclk_205580), .D (n_26), .Q
       (n_4754));
  DFRQX1 \integer_file_reg[13][10] (.C (rc_gclk_205580), .D (n_62), .Q
       (n_5095));
  DFRQX1 \integer_file_reg[13][11] (.C (rc_gclk_205580), .D (n_66), .Q
       (n_5126));
  DFRQX1 \integer_file_reg[13][12] (.C (rc_gclk_205580), .D (n_28), .Q
       (n_5157));
  DFRQX1 \integer_file_reg[13][13] (.C (rc_gclk_205580), .D (n_54), .Q
       (n_5219));
  DFRQX1 \integer_file_reg[13][14] (.C (rc_gclk_205580), .D (n_37), .Q
       (n_5250));
  DFRQX1 \integer_file_reg[13][15] (.C (rc_gclk_205580), .D (n_53), .Q
       (n_5281));
  DFRQX1 \integer_file_reg[13][16] (.C (rc_gclk_205580), .D (n_65), .Q
       (n_5312));
  DFRQX1 \integer_file_reg[13][17] (.C (rc_gclk_205580), .D (n_61), .Q
       (n_5343));
  DFRQX1 \integer_file_reg[13][18] (.C (rc_gclk_205580), .D (n_43), .Q
       (n_5374));
  DFRQX1 \integer_file_reg[13][19] (.C (rc_gclk_205580), .D (n_51), .Q
       (n_5405));
  DFRQX1 \integer_file_reg[13][1] (.C (rc_gclk_205580), .D (n_18), .Q
       (n_4785));
  DFRQX1 \integer_file_reg[13][20] (.C (rc_gclk_205580), .D (n_60), .Q
       (n_5436));
  DFRQX1 \integer_file_reg[13][21] (.C (rc_gclk_205580), .D (n_59), .Q
       (n_5467));
  DFRQX1 \integer_file_reg[13][22] (.C (rc_gclk_205580), .D (n_72), .Q
       (n_5498));
  DFRQX1 \integer_file_reg[13][23] (.C (rc_gclk_205580), .D (n_71), .Q
       (n_4568));
  DFRQX1 \integer_file_reg[13][24] (.C (rc_gclk_205580), .D (n_70), .Q
       (n_4599));
  DFRQX1 \integer_file_reg[13][25] (.C (rc_gclk_205580), .D (n_36), .Q
       (n_4630));
  DFRQX1 \integer_file_reg[13][26] (.C (rc_gclk_205580), .D (n_35), .Q
       (n_4661));
  DFRQX1 \integer_file_reg[13][27] (.C (rc_gclk_205580), .D (n_69), .Q
       (n_4692));
  DFRQX1 \integer_file_reg[13][28] (.C (rc_gclk_205580), .D (n_41), .Q
       (n_4723));
  DFRQX1 \integer_file_reg[13][29] (.C (rc_gclk_205580), .D (n_49), .Q
       (n_4847));
  DFRQX1 \integer_file_reg[13][2] (.C (rc_gclk_205580), .D (n_17), .Q
       (n_4816));
  DFRQX1 \integer_file_reg[13][30] (.C (rc_gclk_205580), .D (n_48), .Q
       (n_5188));
  DFRQX1 \integer_file_reg[13][31] (.C (rc_gclk_205580), .D (n_63), .Q
       (n_5529));
  DFRQX1 \integer_file_reg[13][3] (.C (rc_gclk_205580), .D (n_25), .Q
       (n_4878));
  DFRQX1 \integer_file_reg[13][4] (.C (rc_gclk_205580), .D (n_24), .Q
       (n_4909));
  DFRQX1 \integer_file_reg[13][5] (.C (rc_gclk_205580), .D (n_34), .Q
       (n_4940));
  DFRQX1 \integer_file_reg[13][6] (.C (rc_gclk_205580), .D (n_23), .Q
       (n_4971));
  DFRQX1 \integer_file_reg[13][7] (.C (rc_gclk_205580), .D (n_33), .Q
       (n_5002));
  DFRQX1 \integer_file_reg[13][8] (.C (rc_gclk_205580), .D (n_57), .Q
       (n_5033));
  DFRQX1 \integer_file_reg[13][9] (.C (rc_gclk_205580), .D (n_47), .Q
       (n_5064));
  DFRQX1 \integer_file_reg[14][0] (.C (rc_gclk_205589), .D (n_21), .Q
       (n_4753));
  DFRQX1 \integer_file_reg[14][10] (.C (rc_gclk_205589), .D (n_78), .Q
       (n_5094));
  DFRQX1 \integer_file_reg[14][11] (.C (rc_gclk_205589), .D (n_77), .Q
       (n_5125));
  DFRQX1 \integer_file_reg[14][12] (.C (rc_gclk_205589), .D (n_38), .Q
       (n_5156));
  DFRQX1 \integer_file_reg[14][13] (.C (rc_gclk_205589), .D (n_44), .Q
       (n_5218));
  DFRQX1 \integer_file_reg[14][14] (.C (rc_gclk_205589), .D (n_32), .Q
       (n_5249));
  DFRQX1 \integer_file_reg[14][15] (.C (rc_gclk_205589), .D (n_53), .Q
       (n_5280));
  DFRQX1 \integer_file_reg[14][16] (.C (rc_gclk_205589), .D (n_65), .Q
       (n_5311));
  DFRQX1 \integer_file_reg[14][17] (.C (rc_gclk_205589), .D (n_75), .Q
       (n_5342));
  DFRQX1 \integer_file_reg[14][18] (.C (rc_gclk_205589), .D (n_43), .Q
       (n_5373));
  DFRQX1 \integer_file_reg[14][19] (.C (rc_gclk_205589), .D (n_51), .Q
       (n_5404));
  DFRQX1 \integer_file_reg[14][1] (.C (rc_gclk_205589), .D (n_15), .Q
       (n_4784));
  DFRQX1 \integer_file_reg[14][20] (.C (rc_gclk_205589), .D (n_60), .Q
       (n_5435));
  DFRQX1 \integer_file_reg[14][21] (.C (rc_gclk_205589), .D (n_73), .Q
       (n_5466));
  DFRQX1 \integer_file_reg[14][22] (.C (rc_gclk_205589), .D (n_72), .Q
       (n_5497));
  DFRQX1 \integer_file_reg[14][23] (.C (rc_gclk_205589), .D (n_71), .Q
       (n_4567));
  DFRQX1 \integer_file_reg[14][24] (.C (rc_gclk_205589), .D (n_64), .Q
       (n_4598));
  DFRQX1 \integer_file_reg[14][25] (.C (rc_gclk_205589), .D (n_36), .Q
       (n_4629));
  DFRQX1 \integer_file_reg[14][26] (.C (rc_gclk_205589), .D (n_35), .Q
       (n_4660));
  DFRQX1 \integer_file_reg[14][27] (.C (rc_gclk_205589), .D (n_69), .Q
       (n_4691));
  DFRQX1 \integer_file_reg[14][28] (.C (rc_gclk_205589), .D (n_50), .Q
       (n_4722));
  DFRQX1 \integer_file_reg[14][29] (.C (rc_gclk_205589), .D (n_49), .Q
       (n_4846));
  DFRQX1 \integer_file_reg[14][2] (.C (rc_gclk_205589), .D (n_16), .Q
       (n_4815));
  DFRQX1 \integer_file_reg[14][30] (.C (rc_gclk_205589), .D (n_45), .Q
       (n_5187));
  DFRQX1 \integer_file_reg[14][31] (.C (rc_gclk_205589), .D (n_63), .Q
       (n_5528));
  DFRQX1 \integer_file_reg[14][3] (.C (rc_gclk_205589), .D (n_25), .Q
       (n_4877));
  DFRQX1 \integer_file_reg[14][4] (.C (rc_gclk_205589), .D (n_22), .Q
       (n_4908));
  DFRQX1 \integer_file_reg[14][5] (.C (rc_gclk_205589), .D (n_34), .Q
       (n_4939));
  DFRQX1 \integer_file_reg[14][6] (.C (rc_gclk_205589), .D (n_20), .Q
       (n_4970));
  DFRQX1 \integer_file_reg[14][7] (.C (rc_gclk_205589), .D (n_33), .Q
       (n_5001));
  DFRQX1 \integer_file_reg[14][8] (.C (rc_gclk_205589), .D (n_57), .Q
       (n_5032));
  DFRQX1 \integer_file_reg[14][9] (.C (rc_gclk_205589), .D (n_40), .Q
       (n_5063));
  DFRQX1 \integer_file_reg[15][0] (.C (rc_gclk_205499), .D (n_26), .Q
       (n_4752));
  DFRQX1 \integer_file_reg[15][10] (.C (rc_gclk_205499), .D (n_78), .Q
       (n_5093));
  DFRQX1 \integer_file_reg[15][11] (.C (rc_gclk_205499), .D (n_66), .Q
       (n_5124));
  DFRQX1 \integer_file_reg[15][12] (.C (rc_gclk_205499), .D (n_38), .Q
       (n_5155));
  DFRQX1 \integer_file_reg[15][13] (.C (rc_gclk_205499), .D (n_44), .Q
       (n_5217));
  DFRQX1 \integer_file_reg[15][14] (.C (rc_gclk_205499), .D (n_37), .Q
       (n_5248));
  DFRQX1 \integer_file_reg[15][15] (.C (rc_gclk_205499), .D (n_53), .Q
       (n_5279));
  DFRQX1 \integer_file_reg[15][16] (.C (rc_gclk_205499), .D (n_76), .Q
       (n_5310));
  DFRQX1 \integer_file_reg[15][17] (.C (rc_gclk_205499), .D (n_61), .Q
       (n_5341));
  DFRQX1 \integer_file_reg[15][18] (.C (rc_gclk_205499), .D (n_52), .Q
       (n_5372));
  DFRQX1 \integer_file_reg[15][19] (.C (rc_gclk_205499), .D (n_51), .Q
       (n_5403));
  DFRQX1 \integer_file_reg[15][1] (.C (rc_gclk_205499), .D (n_15), .Q
       (n_4783));
  DFRQX1 \integer_file_reg[15][20] (.C (rc_gclk_205499), .D (n_60), .Q
       (n_5434));
  DFRQX1 \integer_file_reg[15][21] (.C (rc_gclk_205499), .D (n_59), .Q
       (n_5465));
  DFRQX1 \integer_file_reg[15][22] (.C (rc_gclk_205499), .D (n_72), .Q
       (n_5496));
  DFRQX1 \integer_file_reg[15][23] (.C (rc_gclk_205499), .D (n_71), .Q
       (n_4566));
  DFRQX1 \integer_file_reg[15][24] (.C (rc_gclk_205499), .D (n_64), .Q
       (n_4597));
  DFRQX1 \integer_file_reg[15][25] (.C (rc_gclk_205499), .D (n_27), .Q
       (n_4628));
  DFRQX1 \integer_file_reg[15][26] (.C (rc_gclk_205499), .D (n_31), .Q
       (n_4659));
  DFRQX1 \integer_file_reg[15][27] (.C (rc_gclk_205499), .D (n_58), .Q
       (n_4690));
  DFRQX1 \integer_file_reg[15][28] (.C (rc_gclk_205499), .D (n_41), .Q
       (n_4721));
  DFRQX1 \integer_file_reg[15][29] (.C (rc_gclk_205499), .D (n_49), .Q
       (n_4845));
  DFRQX1 \integer_file_reg[15][2] (.C (rc_gclk_205499), .D (n_17), .Q
       (n_4814));
  DFRQX1 \integer_file_reg[15][30] (.C (rc_gclk_205499), .D (n_48), .Q
       (n_5186));
  DFRQX1 \integer_file_reg[15][31] (.C (rc_gclk_205499), .D (n_63), .Q
       (n_5527));
  DFRQX1 \integer_file_reg[15][3] (.C (rc_gclk_205499), .D (n_19), .Q
       (n_4876));
  DFRQX1 \integer_file_reg[15][4] (.C (rc_gclk_205499), .D (n_22), .Q
       (n_4907));
  DFRQX1 \integer_file_reg[15][5] (.C (rc_gclk_205499), .D (n_30), .Q
       (n_4938));
  DFRQX1 \integer_file_reg[15][6] (.C (rc_gclk_205499), .D (n_23), .Q
       (n_4969));
  DFRQX1 \integer_file_reg[15][7] (.C (rc_gclk_205499), .D (n_29), .Q
       (n_5000));
  DFRQX1 \integer_file_reg[15][8] (.C (rc_gclk_205499), .D (n_67), .Q
       (n_5031));
  DFRQX1 \integer_file_reg[15][9] (.C (rc_gclk_205499), .D (n_47), .Q
       (n_5062));
  DFRQX1 \integer_file_reg[16][0] (.C (rc_gclk_205508), .D (n_26), .Q
       (n_4751));
  DFRQX1 \integer_file_reg[16][10] (.C (rc_gclk_205508), .D (n_78), .Q
       (n_5092));
  DFRQX1 \integer_file_reg[16][11] (.C (rc_gclk_205508), .D (n_77), .Q
       (n_5123));
  DFRQX1 \integer_file_reg[16][12] (.C (rc_gclk_205508), .D (n_38), .Q
       (n_5154));
  DFRQX1 \integer_file_reg[16][13] (.C (rc_gclk_205508), .D (n_44), .Q
       (n_5216));
  DFRQX1 \integer_file_reg[16][14] (.C (rc_gclk_205508), .D (n_37), .Q
       (n_5247));
  DFRQX1 \integer_file_reg[16][15] (.C (rc_gclk_205508), .D (n_53), .Q
       (n_5278));
  DFRQX1 \integer_file_reg[16][16] (.C (rc_gclk_205508), .D (n_65), .Q
       (n_5309));
  DFRQX1 \integer_file_reg[16][17] (.C (rc_gclk_205508), .D (n_61), .Q
       (n_5340));
  DFRQX1 \integer_file_reg[16][18] (.C (rc_gclk_205508), .D (n_52), .Q
       (n_5371));
  DFRQX1 \integer_file_reg[16][19] (.C (rc_gclk_205508), .D (n_39), .Q
       (n_5402));
  DFRQX1 \integer_file_reg[16][1] (.C (rc_gclk_205508), .D (n_15), .Q
       (n_4782));
  DFRQX1 \integer_file_reg[16][20] (.C (rc_gclk_205508), .D (n_60), .Q
       (n_5433));
  DFRQX1 \integer_file_reg[16][21] (.C (rc_gclk_205508), .D (n_59), .Q
       (n_5464));
  DFRQX1 \integer_file_reg[16][22] (.C (rc_gclk_205508), .D (n_72), .Q
       (n_5495));
  DFRQX1 \integer_file_reg[16][23] (.C (rc_gclk_205508), .D (n_71), .Q
       (n_4565));
  DFRQX1 \integer_file_reg[16][24] (.C (rc_gclk_205508), .D (n_64), .Q
       (n_4596));
  DFRQX1 \integer_file_reg[16][25] (.C (rc_gclk_205508), .D (n_36), .Q
       (n_4627));
  DFRQX1 \integer_file_reg[16][26] (.C (rc_gclk_205508), .D (n_31), .Q
       (n_4658));
  DFRQX1 \integer_file_reg[16][27] (.C (rc_gclk_205508), .D (n_69), .Q
       (n_4689));
  DFRQX1 \integer_file_reg[16][28] (.C (rc_gclk_205508), .D (n_41), .Q
       (n_4720));
  DFRQX1 \integer_file_reg[16][29] (.C (rc_gclk_205508), .D (n_42), .Q
       (n_4844));
  DFRQX1 \integer_file_reg[16][2] (.C (rc_gclk_205508), .D (n_16), .Q
       (n_4813));
  DFRQX1 \integer_file_reg[16][30] (.C (rc_gclk_205508), .D (n_48), .Q
       (n_5185));
  DFRQX1 \integer_file_reg[16][31] (.C (rc_gclk_205508), .D (n_63), .Q
       (n_5526));
  DFRQX1 \integer_file_reg[16][3] (.C (rc_gclk_205508), .D (n_25), .Q
       (n_4875));
  DFRQX1 \integer_file_reg[16][4] (.C (rc_gclk_205508), .D (n_22), .Q
       (n_4906));
  DFRQX1 \integer_file_reg[16][5] (.C (rc_gclk_205508), .D (n_34), .Q
       (n_4937));
  DFRQX1 \integer_file_reg[16][6] (.C (rc_gclk_205508), .D (n_23), .Q
       (n_4968));
  DFRQX1 \integer_file_reg[16][7] (.C (rc_gclk_205508), .D (n_33), .Q
       (n_4999));
  DFRQX1 \integer_file_reg[16][8] (.C (rc_gclk_205508), .D (n_67), .Q
       (n_5030));
  DFRQX1 \integer_file_reg[16][9] (.C (rc_gclk_205508), .D (n_47), .Q
       (n_5061));
  DFRQX1 \integer_file_reg[17][0] (.C (rc_gclk_205517), .D (n_26), .Q
       (n_4750));
  DFRQX1 \integer_file_reg[17][10] (.C (rc_gclk_205517), .D (n_78), .Q
       (n_5091));
  DFRQX1 \integer_file_reg[17][11] (.C (rc_gclk_205517), .D (n_66), .Q
       (n_5122));
  DFRQX1 \integer_file_reg[17][12] (.C (rc_gclk_205517), .D (n_38), .Q
       (n_5153));
  DFRQX1 \integer_file_reg[17][13] (.C (rc_gclk_205517), .D (n_44), .Q
       (n_5215));
  DFRQX1 \integer_file_reg[17][14] (.C (rc_gclk_205517), .D (n_37), .Q
       (n_5246));
  DFRQX1 \integer_file_reg[17][15] (.C (rc_gclk_205517), .D (n_46), .Q
       (n_5277));
  DFRQX1 \integer_file_reg[17][16] (.C (rc_gclk_205517), .D (n_65), .Q
       (n_5308));
  DFRQX1 \integer_file_reg[17][17] (.C (rc_gclk_205517), .D (n_75), .Q
       (n_5339));
  DFRQX1 \integer_file_reg[17][18] (.C (rc_gclk_205517), .D (n_52), .Q
       (n_5370));
  DFRQX1 \integer_file_reg[17][19] (.C (rc_gclk_205517), .D (n_51), .Q
       (n_5401));
  DFRQX1 \integer_file_reg[17][1] (.C (rc_gclk_205517), .D (n_15), .Q
       (n_4781));
  DFRQX1 \integer_file_reg[17][20] (.C (rc_gclk_205517), .D (n_60), .Q
       (n_5432));
  DFRQX1 \integer_file_reg[17][21] (.C (rc_gclk_205517), .D (n_73), .Q
       (n_5463));
  DFRQX1 \integer_file_reg[17][22] (.C (rc_gclk_205517), .D (n_72), .Q
       (n_5494));
  DFRQX1 \integer_file_reg[17][23] (.C (rc_gclk_205517), .D (n_71), .Q
       (n_4564));
  DFRQX1 \integer_file_reg[17][24] (.C (rc_gclk_205517), .D (n_64), .Q
       (n_4595));
  DFRQX1 \integer_file_reg[17][25] (.C (rc_gclk_205517), .D (n_27), .Q
       (n_4626));
  DFRQX1 \integer_file_reg[17][26] (.C (rc_gclk_205517), .D (n_31), .Q
       (n_4657));
  DFRQX1 \integer_file_reg[17][27] (.C (rc_gclk_205517), .D (n_69), .Q
       (n_4688));
  DFRQX1 \integer_file_reg[17][28] (.C (rc_gclk_205517), .D (n_50), .Q
       (n_4719));
  DFRQX1 \integer_file_reg[17][29] (.C (rc_gclk_205517), .D (n_49), .Q
       (n_4843));
  DFRQX1 \integer_file_reg[17][2] (.C (rc_gclk_205517), .D (n_16), .Q
       (n_4812));
  DFRQX1 \integer_file_reg[17][30] (.C (rc_gclk_205517), .D (n_45), .Q
       (n_5184));
  DFRQX1 \integer_file_reg[17][31] (.C (rc_gclk_205517), .D (n_63), .Q
       (n_5525));
  DFRQX1 \integer_file_reg[17][3] (.C (rc_gclk_205517), .D (n_25), .Q
       (n_4874));
  DFRQX1 \integer_file_reg[17][4] (.C (rc_gclk_205517), .D (n_22), .Q
       (n_4905));
  DFRQX1 \integer_file_reg[17][5] (.C (rc_gclk_205517), .D (n_30), .Q
       (n_4936));
  DFRQX1 \integer_file_reg[17][6] (.C (rc_gclk_205517), .D (n_23), .Q
       (n_4967));
  DFRQX1 \integer_file_reg[17][7] (.C (rc_gclk_205517), .D (n_33), .Q
       (n_4998));
  DFRQX1 \integer_file_reg[17][8] (.C (rc_gclk_205517), .D (n_67), .Q
       (n_5029));
  DFRQX1 \integer_file_reg[17][9] (.C (rc_gclk_205517), .D (n_47), .Q
       (n_5060));
  DFRQX1 \integer_file_reg[18][0] (.C (rc_gclk_205526), .D (n_21), .Q
       (n_4749));
  DFRQX1 \integer_file_reg[18][10] (.C (rc_gclk_205526), .D (n_62), .Q
       (n_5090));
  DFRQX1 \integer_file_reg[18][11] (.C (rc_gclk_205526), .D (n_66), .Q
       (n_5121));
  DFRQX1 \integer_file_reg[18][12] (.C (rc_gclk_205526), .D (n_38), .Q
       (n_5152));
  DFRQX1 \integer_file_reg[18][13] (.C (rc_gclk_205526), .D (n_44), .Q
       (n_5214));
  DFRQX1 \integer_file_reg[18][14] (.C (rc_gclk_205526), .D (n_37), .Q
       (n_5245));
  DFRQX1 \integer_file_reg[18][15] (.C (rc_gclk_205526), .D (n_53), .Q
       (n_5276));
  DFRQX1 \integer_file_reg[18][16] (.C (rc_gclk_205526), .D (n_76), .Q
       (n_5307));
  DFRQX1 \integer_file_reg[18][17] (.C (rc_gclk_205526), .D (n_61), .Q
       (n_5338));
  DFRQX1 \integer_file_reg[18][18] (.C (rc_gclk_205526), .D (n_43), .Q
       (n_5369));
  DFRQX1 \integer_file_reg[18][19] (.C (rc_gclk_205526), .D (n_51), .Q
       (n_5400));
  DFRQX1 \integer_file_reg[18][1] (.C (rc_gclk_205526), .D (n_15), .Q
       (n_4780));
  DFRQX1 \integer_file_reg[18][20] (.C (rc_gclk_205526), .D (n_74), .Q
       (n_5431));
  DFRQX1 \integer_file_reg[18][21] (.C (rc_gclk_205526), .D (n_59), .Q
       (n_5462));
  DFRQX1 \integer_file_reg[18][22] (.C (rc_gclk_205526), .D (n_72), .Q
       (n_5493));
  DFRQX1 \integer_file_reg[18][23] (.C (rc_gclk_205526), .D (n_71), .Q
       (n_4563));
  DFRQX1 \integer_file_reg[18][24] (.C (rc_gclk_205526), .D (n_64), .Q
       (n_4594));
  DFRQX1 \integer_file_reg[18][25] (.C (rc_gclk_205526), .D (n_27), .Q
       (n_4625));
  DFRQX1 \integer_file_reg[18][26] (.C (rc_gclk_205526), .D (n_35), .Q
       (n_4656));
  DFRQX1 \integer_file_reg[18][27] (.C (rc_gclk_205526), .D (n_69), .Q
       (n_4687));
  DFRQX1 \integer_file_reg[18][28] (.C (rc_gclk_205526), .D (n_50), .Q
       (n_4718));
  DFRQX1 \integer_file_reg[18][29] (.C (rc_gclk_205526), .D (n_42), .Q
       (n_4842));
  DFRQX1 \integer_file_reg[18][2] (.C (rc_gclk_205526), .D (n_17), .Q
       (n_4811));
  DFRQX1 \integer_file_reg[18][30] (.C (rc_gclk_205526), .D (n_48), .Q
       (n_5183));
  DFRQX1 \integer_file_reg[18][31] (.C (rc_gclk_205526), .D (n_63), .Q
       (n_5524));
  DFRQX1 \integer_file_reg[18][3] (.C (rc_gclk_205526), .D (n_19), .Q
       (n_4873));
  DFRQX1 \integer_file_reg[18][4] (.C (rc_gclk_205526), .D (n_24), .Q
       (n_4904));
  DFRQX1 \integer_file_reg[18][5] (.C (rc_gclk_205526), .D (n_30), .Q
       (n_4935));
  DFRQX1 \integer_file_reg[18][6] (.C (rc_gclk_205526), .D (n_23), .Q
       (n_4966));
  DFRQX1 \integer_file_reg[18][7] (.C (rc_gclk_205526), .D (n_33), .Q
       (n_4997));
  DFRQX1 \integer_file_reg[18][8] (.C (rc_gclk_205526), .D (n_67), .Q
       (n_5028));
  DFRQX1 \integer_file_reg[18][9] (.C (rc_gclk_205526), .D (n_47), .Q
       (n_5059));
  DFRQX1 \integer_file_reg[19][0] (.C (rc_gclk_205538), .D (n_21), .Q
       (n_4748));
  DFRQX1 \integer_file_reg[19][10] (.C (rc_gclk_205538), .D (n_78), .Q
       (n_5089));
  DFRQX1 \integer_file_reg[19][11] (.C (rc_gclk_205538), .D (n_66), .Q
       (n_5120));
  DFRQX1 \integer_file_reg[19][12] (.C (rc_gclk_205538), .D (n_28), .Q
       (n_5151));
  DFRQX1 \integer_file_reg[19][13] (.C (rc_gclk_205538), .D (n_44), .Q
       (n_5213));
  DFRQX1 \integer_file_reg[19][14] (.C (rc_gclk_205538), .D (n_32), .Q
       (n_5244));
  DFRQX1 \integer_file_reg[19][15] (.C (rc_gclk_205538), .D (n_53), .Q
       (n_5275));
  DFRQX1 \integer_file_reg[19][16] (.C (rc_gclk_205538), .D (n_65), .Q
       (n_5306));
  DFRQX1 \integer_file_reg[19][17] (.C (rc_gclk_205538), .D (n_61), .Q
       (n_5337));
  DFRQX1 \integer_file_reg[19][18] (.C (rc_gclk_205538), .D (n_43), .Q
       (n_5368));
  DFRQX1 \integer_file_reg[19][19] (.C (rc_gclk_205538), .D (n_39), .Q
       (n_5399));
  DFRQX1 \integer_file_reg[19][1] (.C (rc_gclk_205538), .D (n_15), .Q
       (n_4779));
  DFRQX1 \integer_file_reg[19][20] (.C (rc_gclk_205538), .D (n_74), .Q
       (n_5430));
  DFRQX1 \integer_file_reg[19][21] (.C (rc_gclk_205538), .D (n_59), .Q
       (n_5461));
  DFRQX1 \integer_file_reg[19][22] (.C (rc_gclk_205538), .D (n_56), .Q
       (n_5492));
  DFRQX1 \integer_file_reg[19][23] (.C (rc_gclk_205538), .D (n_71), .Q
       (n_4562));
  DFRQX1 \integer_file_reg[19][24] (.C (rc_gclk_205538), .D (n_64), .Q
       (n_4593));
  DFRQX1 \integer_file_reg[19][25] (.C (rc_gclk_205538), .D (n_27), .Q
       (n_4624));
  DFRQX1 \integer_file_reg[19][26] (.C (rc_gclk_205538), .D (n_31), .Q
       (n_4655));
  DFRQX1 \integer_file_reg[19][27] (.C (rc_gclk_205538), .D (n_69), .Q
       (n_4686));
  DFRQX1 \integer_file_reg[19][28] (.C (rc_gclk_205538), .D (n_41), .Q
       (n_4717));
  DFRQX1 \integer_file_reg[19][29] (.C (rc_gclk_205538), .D (n_42), .Q
       (n_4841));
  DFRQX1 \integer_file_reg[19][2] (.C (rc_gclk_205538), .D (n_17), .Q
       (n_4810));
  DFRQX1 \integer_file_reg[19][30] (.C (rc_gclk_205538), .D (n_48), .Q
       (n_5182));
  DFRQX1 \integer_file_reg[19][31] (.C (rc_gclk_205538), .D (n_63), .Q
       (n_5523));
  DFRQX1 \integer_file_reg[19][3] (.C (rc_gclk_205538), .D (n_19), .Q
       (n_4872));
  DFRQX1 \integer_file_reg[19][4] (.C (rc_gclk_205538), .D (n_22), .Q
       (n_4903));
  DFRQX1 \integer_file_reg[19][5] (.C (rc_gclk_205538), .D (n_30), .Q
       (n_4934));
  DFRQX1 \integer_file_reg[19][6] (.C (rc_gclk_205538), .D (n_23), .Q
       (n_4965));
  DFRQX1 \integer_file_reg[19][7] (.C (rc_gclk_205538), .D (n_29), .Q
       (n_4996));
  DFRQX1 \integer_file_reg[19][8] (.C (rc_gclk_205538), .D (n_67), .Q
       (n_5027));
  DFRQX1 \integer_file_reg[19][9] (.C (rc_gclk_205538), .D (n_47), .Q
       (n_5058));
  DFRQX1 \integer_file_reg[1][0] (.C (rc_gclk_205547), .D (n_21), .Q
       (n_4766));
  DFRQX1 \integer_file_reg[1][10] (.C (rc_gclk_205547), .D (n_78), .Q
       (n_5107));
  DFRQX1 \integer_file_reg[1][11] (.C (rc_gclk_205547), .D (n_66), .Q
       (n_5138));
  DFRQX1 \integer_file_reg[1][12] (.C (rc_gclk_205547), .D (n_28), .Q
       (n_5169));
  DFRQX1 \integer_file_reg[1][13] (.C (rc_gclk_205547), .D (n_44), .Q
       (n_5231));
  DFRQX1 \integer_file_reg[1][14] (.C (rc_gclk_205547), .D (n_32), .Q
       (n_5262));
  DFRQX1 \integer_file_reg[1][15] (.C (rc_gclk_205547), .D (n_46), .Q
       (n_5293));
  DFRQX1 \integer_file_reg[1][16] (.C (rc_gclk_205547), .D (n_65), .Q
       (n_5324));
  DFRQX1 \integer_file_reg[1][17] (.C (rc_gclk_205547), .D (n_61), .Q
       (n_5355));
  DFRQX1 \integer_file_reg[1][18] (.C (rc_gclk_205547), .D (n_52), .Q
       (n_5386));
  DFRQX1 \integer_file_reg[1][19] (.C (rc_gclk_205547), .D (n_51), .Q
       (n_5417));
  DFRQX1 \integer_file_reg[1][1] (.C (rc_gclk_205547), .D (n_15), .Q
       (n_4797));
  DFRQX1 \integer_file_reg[1][20] (.C (rc_gclk_205547), .D (n_60), .Q
       (n_5448));
  DFRQX1 \integer_file_reg[1][21] (.C (rc_gclk_205547), .D (n_73), .Q
       (n_5479));
  DFRQX1 \integer_file_reg[1][22] (.C (rc_gclk_205547), .D (n_72), .Q
       (n_5510));
  DFRQX1 \integer_file_reg[1][23] (.C (rc_gclk_205547), .D (n_71), .Q
       (n_4580));
  DFRQX1 \integer_file_reg[1][24] (.C (rc_gclk_205547), .D (n_64), .Q
       (n_4611));
  DFRQX1 \integer_file_reg[1][25] (.C (rc_gclk_205547), .D (n_36), .Q
       (n_4642));
  DFRQX1 \integer_file_reg[1][26] (.C (rc_gclk_205547), .D (n_31), .Q
       (n_4673));
  DFRQX1 \integer_file_reg[1][27] (.C (rc_gclk_205547), .D (n_69), .Q
       (n_4704));
  DFRQX1 \integer_file_reg[1][28] (.C (rc_gclk_205547), .D (n_41), .Q
       (n_4735));
  DFRQX1 \integer_file_reg[1][29] (.C (rc_gclk_205547), .D (n_42), .Q
       (n_4859));
  DFRQX1 \integer_file_reg[1][2] (.C (rc_gclk_205547), .D (n_16), .Q
       (n_4828));
  DFRQX1 \integer_file_reg[1][30] (.C (rc_gclk_205547), .D (n_48), .Q
       (n_5200));
  DFRQX1 \integer_file_reg[1][31] (.C (rc_gclk_205547), .D (n_63), .Q
       (n_5541));
  DFRQX1 \integer_file_reg[1][3] (.C (rc_gclk_205547), .D (n_25), .Q
       (n_4890));
  DFRQX1 \integer_file_reg[1][4] (.C (rc_gclk_205547), .D (n_22), .Q
       (n_4921));
  DFRQX1 \integer_file_reg[1][5] (.C (rc_gclk_205547), .D (n_34), .Q
       (n_4952));
  DFRQX1 \integer_file_reg[1][6] (.C (rc_gclk_205547), .D (n_23), .Q
       (n_4983));
  DFRQX1 \integer_file_reg[1][7] (.C (rc_gclk_205547), .D (n_29), .Q
       (n_5014));
  DFRQX1 \integer_file_reg[1][8] (.C (rc_gclk_205547), .D (n_57), .Q
       (n_5045));
  DFRQX1 \integer_file_reg[1][9] (.C (rc_gclk_205547), .D (n_47), .Q
       (n_5076));
  DFRQX1 \integer_file_reg[20][0] (.C (rc_gclk_205550), .D (n_26), .Q
       (n_4747));
  DFRQX1 \integer_file_reg[20][10] (.C (rc_gclk_205550), .D (n_78), .Q
       (n_5088));
  DFRQX1 \integer_file_reg[20][11] (.C (rc_gclk_205550), .D (n_66), .Q
       (n_5119));
  DFRQX1 \integer_file_reg[20][12] (.C (rc_gclk_205550), .D (n_38), .Q
       (n_5150));
  DFRQX1 \integer_file_reg[20][13] (.C (rc_gclk_205550), .D (n_54), .Q
       (n_5212));
  DFRQX1 \integer_file_reg[20][14] (.C (rc_gclk_205550), .D (n_32), .Q
       (n_5243));
  DFRQX1 \integer_file_reg[20][15] (.C (rc_gclk_205550), .D (n_53), .Q
       (n_5274));
  DFRQX1 \integer_file_reg[20][16] (.C (rc_gclk_205550), .D (n_65), .Q
       (n_5305));
  DFRQX1 \integer_file_reg[20][17] (.C (rc_gclk_205550), .D (n_75), .Q
       (n_5336));
  DFRQX1 \integer_file_reg[20][18] (.C (rc_gclk_205550), .D (n_43), .Q
       (n_5367));
  DFRQX1 \integer_file_reg[20][19] (.C (rc_gclk_205550), .D (n_51), .Q
       (n_5398));
  DFRQX1 \integer_file_reg[20][1] (.C (rc_gclk_205550), .D (n_15), .Q
       (n_4778));
  DFRQX1 \integer_file_reg[20][20] (.C (rc_gclk_205550), .D (n_60), .Q
       (n_5429));
  DFRQX1 \integer_file_reg[20][21] (.C (rc_gclk_205550), .D (n_73), .Q
       (n_5460));
  DFRQX1 \integer_file_reg[20][22] (.C (rc_gclk_205550), .D (n_72), .Q
       (n_5491));
  DFRQX1 \integer_file_reg[20][23] (.C (rc_gclk_205550), .D (n_71), .Q
       (n_4561));
  DFRQX1 \integer_file_reg[20][24] (.C (rc_gclk_205550), .D (n_64), .Q
       (n_4592));
  DFRQX1 \integer_file_reg[20][25] (.C (rc_gclk_205550), .D (n_27), .Q
       (n_4623));
  DFRQX1 \integer_file_reg[20][26] (.C (rc_gclk_205550), .D (n_31), .Q
       (n_4654));
  DFRQX1 \integer_file_reg[20][27] (.C (rc_gclk_205550), .D (n_69), .Q
       (n_4685));
  DFRQX1 \integer_file_reg[20][28] (.C (rc_gclk_205550), .D (n_50), .Q
       (n_4716));
  DFRQX1 \integer_file_reg[20][29] (.C (rc_gclk_205550), .D (n_49), .Q
       (n_4840));
  DFRQX1 \integer_file_reg[20][2] (.C (rc_gclk_205550), .D (n_17), .Q
       (n_4809));
  DFRQX1 \integer_file_reg[20][30] (.C (rc_gclk_205550), .D (n_45), .Q
       (n_5181));
  DFRQX1 \integer_file_reg[20][31] (.C (rc_gclk_205550), .D (n_63), .Q
       (n_5522));
  DFRQX1 \integer_file_reg[20][3] (.C (rc_gclk_205550), .D (n_25), .Q
       (n_4871));
  DFRQX1 \integer_file_reg[20][4] (.C (rc_gclk_205550), .D (n_22), .Q
       (n_4902));
  DFRQX1 \integer_file_reg[20][5] (.C (rc_gclk_205550), .D (n_34), .Q
       (n_4933));
  DFRQX1 \integer_file_reg[20][6] (.C (rc_gclk_205550), .D (n_23), .Q
       (n_4964));
  DFRQX1 \integer_file_reg[20][7] (.C (rc_gclk_205550), .D (n_33), .Q
       (n_4995));
  DFRQX1 \integer_file_reg[20][8] (.C (rc_gclk_205550), .D (n_67), .Q
       (n_5026));
  DFRQX1 \integer_file_reg[20][9] (.C (rc_gclk_205550), .D (n_47), .Q
       (n_5057));
  DFRQX1 \integer_file_reg[21][0] (.C (rc_gclk_205553), .D (n_21), .Q
       (n_4746));
  DFRQX1 \integer_file_reg[21][10] (.C (rc_gclk_205553), .D (n_78), .Q
       (n_5087));
  DFRQX1 \integer_file_reg[21][11] (.C (rc_gclk_205553), .D (n_77), .Q
       (n_5118));
  DFRQX1 \integer_file_reg[21][12] (.C (rc_gclk_205553), .D (n_38), .Q
       (n_5149));
  DFRQX1 \integer_file_reg[21][13] (.C (rc_gclk_205553), .D (n_54), .Q
       (n_5211));
  DFRQX1 \integer_file_reg[21][14] (.C (rc_gclk_205553), .D (n_37), .Q
       (n_5242));
  DFRQX1 \integer_file_reg[21][15] (.C (rc_gclk_205553), .D (n_53), .Q
       (n_5273));
  DFRQX1 \integer_file_reg[21][16] (.C (rc_gclk_205553), .D (n_65), .Q
       (n_5304));
  DFRQX1 \integer_file_reg[21][17] (.C (rc_gclk_205553), .D (n_61), .Q
       (n_5335));
  DFRQX1 \integer_file_reg[21][18] (.C (rc_gclk_205553), .D (n_43), .Q
       (n_5366));
  DFRQX1 \integer_file_reg[21][19] (.C (rc_gclk_205553), .D (n_51), .Q
       (n_5397));
  DFRQX1 \integer_file_reg[21][1] (.C (rc_gclk_205553), .D (n_15), .Q
       (n_4777));
  DFRQX1 \integer_file_reg[21][20] (.C (rc_gclk_205553), .D (n_74), .Q
       (n_5428));
  DFRQX1 \integer_file_reg[21][21] (.C (rc_gclk_205553), .D (n_73), .Q
       (n_5459));
  DFRQX1 \integer_file_reg[21][22] (.C (rc_gclk_205553), .D (n_72), .Q
       (n_5490));
  DFRQX1 \integer_file_reg[21][23] (.C (rc_gclk_205553), .D (n_71), .Q
       (n_4560));
  DFRQX1 \integer_file_reg[21][24] (.C (rc_gclk_205553), .D (n_64), .Q
       (n_4591));
  DFRQX1 \integer_file_reg[21][25] (.C (rc_gclk_205553), .D (n_36), .Q
       (n_4622));
  DFRQX1 \integer_file_reg[21][26] (.C (rc_gclk_205553), .D (n_31), .Q
       (n_4653));
  DFRQX1 \integer_file_reg[21][27] (.C (rc_gclk_205553), .D (n_69), .Q
       (n_4684));
  DFRQX1 \integer_file_reg[21][28] (.C (rc_gclk_205553), .D (n_50), .Q
       (n_4715));
  DFRQX1 \integer_file_reg[21][29] (.C (rc_gclk_205553), .D (n_42), .Q
       (n_4839));
  DFRQX1 \integer_file_reg[21][2] (.C (rc_gclk_205553), .D (n_17), .Q
       (n_4808));
  DFRQX1 \integer_file_reg[21][30] (.C (rc_gclk_205553), .D (n_48), .Q
       (n_5180));
  DFRQX1 \integer_file_reg[21][31] (.C (rc_gclk_205553), .D (n_63), .Q
       (n_5521));
  DFRQX1 \integer_file_reg[21][3] (.C (rc_gclk_205553), .D (n_25), .Q
       (n_4870));
  DFRQX1 \integer_file_reg[21][4] (.C (rc_gclk_205553), .D (n_22), .Q
       (n_4901));
  DFRQX1 \integer_file_reg[21][5] (.C (rc_gclk_205553), .D (n_34), .Q
       (n_4932));
  DFRQX1 \integer_file_reg[21][6] (.C (rc_gclk_205553), .D (n_20), .Q
       (n_4963));
  DFRQX1 \integer_file_reg[21][7] (.C (rc_gclk_205553), .D (n_33), .Q
       (n_4994));
  DFRQX1 \integer_file_reg[21][8] (.C (rc_gclk_205553), .D (n_67), .Q
       (n_5025));
  DFRQX1 \integer_file_reg[21][9] (.C (rc_gclk_205553), .D (n_47), .Q
       (n_5056));
  DFRQX1 \integer_file_reg[22][0] (.C (rc_gclk_205562), .D (n_26), .Q
       (n_4745));
  DFRQX1 \integer_file_reg[22][10] (.C (rc_gclk_205562), .D (n_62), .Q
       (n_5086));
  DFRQX1 \integer_file_reg[22][11] (.C (rc_gclk_205562), .D (n_66), .Q
       (n_5117));
  DFRQX1 \integer_file_reg[22][12] (.C (rc_gclk_205562), .D (n_38), .Q
       (n_5148));
  DFRQX1 \integer_file_reg[22][13] (.C (rc_gclk_205562), .D (n_54), .Q
       (n_5210));
  DFRQX1 \integer_file_reg[22][14] (.C (rc_gclk_205562), .D (n_37), .Q
       (n_5241));
  DFRQX1 \integer_file_reg[22][15] (.C (rc_gclk_205562), .D (n_53), .Q
       (n_5272));
  DFRQX1 \integer_file_reg[22][16] (.C (rc_gclk_205562), .D (n_76), .Q
       (n_5303));
  DFRQX1 \integer_file_reg[22][17] (.C (rc_gclk_205562), .D (n_61), .Q
       (n_5334));
  DFRQX1 \integer_file_reg[22][18] (.C (rc_gclk_205562), .D (n_43), .Q
       (n_5365));
  DFRQX1 \integer_file_reg[22][19] (.C (rc_gclk_205562), .D (n_39), .Q
       (n_5396));
  DFRQX1 \integer_file_reg[22][1] (.C (rc_gclk_205562), .D (n_15), .Q
       (n_4776));
  DFRQX1 \integer_file_reg[22][20] (.C (rc_gclk_205562), .D (n_60), .Q
       (n_5427));
  DFRQX1 \integer_file_reg[22][21] (.C (rc_gclk_205562), .D (n_73), .Q
       (n_5458));
  DFRQX1 \integer_file_reg[22][22] (.C (rc_gclk_205562), .D (n_72), .Q
       (n_5489));
  DFRQX1 \integer_file_reg[22][23] (.C (rc_gclk_205562), .D (n_71), .Q
       (n_4559));
  DFRQX1 \integer_file_reg[22][24] (.C (rc_gclk_205562), .D (n_64), .Q
       (n_4590));
  DFRQX1 \integer_file_reg[22][25] (.C (rc_gclk_205562), .D (n_36), .Q
       (n_4621));
  DFRQX1 \integer_file_reg[22][26] (.C (rc_gclk_205562), .D (n_31), .Q
       (n_4652));
  DFRQX1 \integer_file_reg[22][27] (.C (rc_gclk_205562), .D (n_69), .Q
       (n_4683));
  DFRQX1 \integer_file_reg[22][28] (.C (rc_gclk_205562), .D (n_50), .Q
       (n_4714));
  DFRQX1 \integer_file_reg[22][29] (.C (rc_gclk_205562), .D (n_42), .Q
       (n_4838));
  DFRQX1 \integer_file_reg[22][2] (.C (rc_gclk_205562), .D (n_17), .Q
       (n_4807));
  DFRQX1 \integer_file_reg[22][30] (.C (rc_gclk_205562), .D (n_45), .Q
       (n_5179));
  DFRQX1 \integer_file_reg[22][31] (.C (rc_gclk_205562), .D (n_63), .Q
       (n_5520));
  DFRQX1 \integer_file_reg[22][3] (.C (rc_gclk_205562), .D (n_25), .Q
       (n_4869));
  DFRQX1 \integer_file_reg[22][4] (.C (rc_gclk_205562), .D (n_22), .Q
       (n_4900));
  DFRQX1 \integer_file_reg[22][5] (.C (rc_gclk_205562), .D (n_34), .Q
       (n_4931));
  DFRQX1 \integer_file_reg[22][6] (.C (rc_gclk_205562), .D (n_20), .Q
       (n_4962));
  DFRQX1 \integer_file_reg[22][7] (.C (rc_gclk_205562), .D (n_33), .Q
       (n_4993));
  DFRQX1 \integer_file_reg[22][8] (.C (rc_gclk_205562), .D (n_67), .Q
       (n_5024));
  DFRQX1 \integer_file_reg[22][9] (.C (rc_gclk_205562), .D (n_47), .Q
       (n_5055));
  DFRQX1 \integer_file_reg[23][0] (.C (rc_gclk_205565), .D (n_21), .Q
       (n_4744));
  DFRQX1 \integer_file_reg[23][10] (.C (rc_gclk_205565), .D (n_62), .Q
       (n_5085));
  DFRQX1 \integer_file_reg[23][11] (.C (rc_gclk_205565), .D (n_77), .Q
       (n_5116));
  DFRQX1 \integer_file_reg[23][12] (.C (rc_gclk_205565), .D (n_38), .Q
       (n_5147));
  DFRQX1 \integer_file_reg[23][13] (.C (rc_gclk_205565), .D (n_54), .Q
       (n_5209));
  DFRQX1 \integer_file_reg[23][14] (.C (rc_gclk_205565), .D (n_32), .Q
       (n_5240));
  DFRQX1 \integer_file_reg[23][15] (.C (rc_gclk_205565), .D (n_53), .Q
       (n_5271));
  DFRQX1 \integer_file_reg[23][16] (.C (rc_gclk_205565), .D (n_65), .Q
       (n_5302));
  DFRQX1 \integer_file_reg[23][17] (.C (rc_gclk_205565), .D (n_61), .Q
       (n_5333));
  DFRQX1 \integer_file_reg[23][18] (.C (rc_gclk_205565), .D (n_52), .Q
       (n_5364));
  DFRQX1 \integer_file_reg[23][19] (.C (rc_gclk_205565), .D (n_39), .Q
       (n_5395));
  DFRQX1 \integer_file_reg[23][1] (.C (rc_gclk_205565), .D (n_15), .Q
       (n_4775));
  DFRQX1 \integer_file_reg[23][20] (.C (rc_gclk_205565), .D (n_60), .Q
       (n_5426));
  DFRQX1 \integer_file_reg[23][21] (.C (rc_gclk_205565), .D (n_73), .Q
       (n_5457));
  DFRQX1 \integer_file_reg[23][22] (.C (rc_gclk_205565), .D (n_72), .Q
       (n_5488));
  DFRQX1 \integer_file_reg[23][23] (.C (rc_gclk_205565), .D (n_71), .Q
       (n_4558));
  DFRQX1 \integer_file_reg[23][24] (.C (rc_gclk_205565), .D (n_64), .Q
       (n_4589));
  DFRQX1 \integer_file_reg[23][25] (.C (rc_gclk_205565), .D (n_36), .Q
       (n_4620));
  DFRQX1 \integer_file_reg[23][26] (.C (rc_gclk_205565), .D (n_31), .Q
       (n_4651));
  DFRQX1 \integer_file_reg[23][27] (.C (rc_gclk_205565), .D (n_69), .Q
       (n_4682));
  DFRQX1 \integer_file_reg[23][28] (.C (rc_gclk_205565), .D (n_50), .Q
       (n_4713));
  DFRQX1 \integer_file_reg[23][29] (.C (rc_gclk_205565), .D (n_49), .Q
       (n_4837));
  DFRQX1 \integer_file_reg[23][2] (.C (rc_gclk_205565), .D (n_17), .Q
       (n_4806));
  DFRQX1 \integer_file_reg[23][30] (.C (rc_gclk_205565), .D (n_45), .Q
       (n_5178));
  DFRQX1 \integer_file_reg[23][31] (.C (rc_gclk_205565), .D (n_63), .Q
       (n_5519));
  DFRQX1 \integer_file_reg[23][3] (.C (rc_gclk_205565), .D (n_19), .Q
       (n_4868));
  DFRQX1 \integer_file_reg[23][4] (.C (rc_gclk_205565), .D (n_24), .Q
       (n_4899));
  DFRQX1 \integer_file_reg[23][5] (.C (rc_gclk_205565), .D (n_34), .Q
       (n_4930));
  DFRQX1 \integer_file_reg[23][6] (.C (rc_gclk_205565), .D (n_23), .Q
       (n_4961));
  DFRQX1 \integer_file_reg[23][7] (.C (rc_gclk_205565), .D (n_29), .Q
       (n_4992));
  DFRQX1 \integer_file_reg[23][8] (.C (rc_gclk_205565), .D (n_57), .Q
       (n_5023));
  DFRQX1 \integer_file_reg[23][9] (.C (rc_gclk_205565), .D (n_47), .Q
       (n_5054));
  DFRQX1 \integer_file_reg[24][0] (.C (rc_gclk_205571), .D (n_26), .Q
       (n_4743));
  DFRQX1 \integer_file_reg[24][10] (.C (rc_gclk_205571), .D (n_78), .Q
       (n_5084));
  DFRQX1 \integer_file_reg[24][11] (.C (rc_gclk_205571), .D (n_66), .Q
       (n_5115));
  DFRQX1 \integer_file_reg[24][12] (.C (rc_gclk_205571), .D (n_38), .Q
       (n_5146));
  DFRQX1 \integer_file_reg[24][13] (.C (rc_gclk_205571), .D (n_54), .Q
       (n_5208));
  DFRQX1 \integer_file_reg[24][14] (.C (rc_gclk_205571), .D (n_37), .Q
       (n_5239));
  DFRQX1 \integer_file_reg[24][15] (.C (rc_gclk_205571), .D (n_53), .Q
       (n_5270));
  DFRQX1 \integer_file_reg[24][16] (.C (rc_gclk_205571), .D (n_65), .Q
       (n_5301));
  DFRQX1 \integer_file_reg[24][17] (.C (rc_gclk_205571), .D (n_75), .Q
       (n_5332));
  DFRQX1 \integer_file_reg[24][18] (.C (rc_gclk_205571), .D (n_43), .Q
       (n_5363));
  DFRQX1 \integer_file_reg[24][19] (.C (rc_gclk_205571), .D (n_51), .Q
       (n_5394));
  DFRQX1 \integer_file_reg[24][1] (.C (rc_gclk_205571), .D (n_15), .Q
       (n_4774));
  DFRQX1 \integer_file_reg[24][20] (.C (rc_gclk_205571), .D (n_74), .Q
       (n_5425));
  DFRQX1 \integer_file_reg[24][21] (.C (rc_gclk_205571), .D (n_59), .Q
       (n_5456));
  DFRQX1 \integer_file_reg[24][22] (.C (rc_gclk_205571), .D (n_72), .Q
       (n_5487));
  DFRQX1 \integer_file_reg[24][23] (.C (rc_gclk_205571), .D (n_55), .Q
       (n_4557));
  DFRQX1 \integer_file_reg[24][24] (.C (rc_gclk_205571), .D (n_70), .Q
       (n_4588));
  DFRQX1 \integer_file_reg[24][25] (.C (rc_gclk_205571), .D (n_27), .Q
       (n_4619));
  DFRQX1 \integer_file_reg[24][26] (.C (rc_gclk_205571), .D (n_31), .Q
       (n_4650));
  DFRQX1 \integer_file_reg[24][27] (.C (rc_gclk_205571), .D (n_69), .Q
       (n_4681));
  DFRQX1 \integer_file_reg[24][28] (.C (rc_gclk_205571), .D (n_41), .Q
       (n_4712));
  DFRQX1 \integer_file_reg[24][29] (.C (rc_gclk_205571), .D (n_49), .Q
       (n_4836));
  DFRQX1 \integer_file_reg[24][2] (.C (rc_gclk_205571), .D (n_17), .Q
       (n_4805));
  DFRQX1 \integer_file_reg[24][30] (.C (rc_gclk_205571), .D (n_48), .Q
       (n_5177));
  DFRQX1 \integer_file_reg[24][31] (.C (rc_gclk_205571), .D (n_63), .Q
       (n_5518));
  DFRQX1 \integer_file_reg[24][3] (.C (rc_gclk_205571), .D (n_25), .Q
       (n_4867));
  DFRQX1 \integer_file_reg[24][4] (.C (rc_gclk_205571), .D (n_22), .Q
       (n_4898));
  DFRQX1 \integer_file_reg[24][5] (.C (rc_gclk_205571), .D (n_34), .Q
       (n_4929));
  DFRQX1 \integer_file_reg[24][6] (.C (rc_gclk_205571), .D (n_23), .Q
       (n_4960));
  DFRQX1 \integer_file_reg[24][7] (.C (rc_gclk_205571), .D (n_33), .Q
       (n_4991));
  DFRQX1 \integer_file_reg[24][8] (.C (rc_gclk_205571), .D (n_67), .Q
       (n_5022));
  DFRQX1 \integer_file_reg[24][9] (.C (rc_gclk_205571), .D (n_47), .Q
       (n_5053));
  DFRQX1 \integer_file_reg[25][0] (.C (rc_gclk_205574), .D (n_26), .Q
       (n_4742));
  DFRQX1 \integer_file_reg[25][10] (.C (rc_gclk_205574), .D (n_62), .Q
       (n_5083));
  DFRQX1 \integer_file_reg[25][11] (.C (rc_gclk_205574), .D (n_66), .Q
       (n_5114));
  DFRQX1 \integer_file_reg[25][12] (.C (rc_gclk_205574), .D (n_28), .Q
       (n_5145));
  DFRQX1 \integer_file_reg[25][13] (.C (rc_gclk_205574), .D (n_44), .Q
       (n_5207));
  DFRQX1 \integer_file_reg[25][14] (.C (rc_gclk_205574), .D (n_37), .Q
       (n_5238));
  DFRQX1 \integer_file_reg[25][15] (.C (rc_gclk_205574), .D (n_53), .Q
       (n_5269));
  DFRQX1 \integer_file_reg[25][16] (.C (rc_gclk_205574), .D (n_65), .Q
       (n_5300));
  DFRQX1 \integer_file_reg[25][17] (.C (rc_gclk_205574), .D (n_61), .Q
       (n_5331));
  DFRQX1 \integer_file_reg[25][18] (.C (rc_gclk_205574), .D (n_43), .Q
       (n_5362));
  DFRQX1 \integer_file_reg[25][19] (.C (rc_gclk_205574), .D (n_51), .Q
       (n_5393));
  DFRQX1 \integer_file_reg[25][1] (.C (rc_gclk_205574), .D (n_15), .Q
       (n_4773));
  DFRQX1 \integer_file_reg[25][20] (.C (rc_gclk_205574), .D (n_74), .Q
       (n_5424));
  DFRQX1 \integer_file_reg[25][21] (.C (rc_gclk_205574), .D (n_73), .Q
       (n_5455));
  DFRQX1 \integer_file_reg[25][22] (.C (rc_gclk_205574), .D (n_72), .Q
       (n_5486));
  DFRQX1 \integer_file_reg[25][23] (.C (rc_gclk_205574), .D (n_71), .Q
       (n_4556));
  DFRQX1 \integer_file_reg[25][24] (.C (rc_gclk_205574), .D (n_70), .Q
       (n_4587));
  DFRQX1 \integer_file_reg[25][25] (.C (rc_gclk_205574), .D (n_36), .Q
       (n_4618));
  DFRQX1 \integer_file_reg[25][26] (.C (rc_gclk_205574), .D (n_31), .Q
       (n_4649));
  DFRQX1 \integer_file_reg[25][27] (.C (rc_gclk_205574), .D (n_69), .Q
       (n_4680));
  DFRQX1 \integer_file_reg[25][28] (.C (rc_gclk_205574), .D (n_41), .Q
       (n_4711));
  DFRQX1 \integer_file_reg[25][29] (.C (rc_gclk_205574), .D (n_42), .Q
       (n_4835));
  DFRQX1 \integer_file_reg[25][2] (.C (rc_gclk_205574), .D (n_16), .Q
       (n_4804));
  DFRQX1 \integer_file_reg[25][30] (.C (rc_gclk_205574), .D (n_45), .Q
       (n_5176));
  DFRQX1 \integer_file_reg[25][31] (.C (rc_gclk_205574), .D (n_63), .Q
       (n_5517));
  DFRQX1 \integer_file_reg[25][3] (.C (rc_gclk_205574), .D (n_25), .Q
       (n_4866));
  DFRQX1 \integer_file_reg[25][4] (.C (rc_gclk_205574), .D (n_24), .Q
       (n_4897));
  DFRQX1 \integer_file_reg[25][5] (.C (rc_gclk_205574), .D (n_34), .Q
       (n_4928));
  DFRQX1 \integer_file_reg[25][6] (.C (rc_gclk_205574), .D (n_23), .Q
       (n_4959));
  DFRQX1 \integer_file_reg[25][7] (.C (rc_gclk_205574), .D (n_33), .Q
       (n_4990));
  DFRQX1 \integer_file_reg[25][8] (.C (rc_gclk_205574), .D (n_57), .Q
       (n_5021));
  DFRQX1 \integer_file_reg[25][9] (.C (rc_gclk_205574), .D (n_40), .Q
       (n_5052));
  DFRQX1 \integer_file_reg[26][0] (.C (rc_gclk_205583), .D (n_21), .Q
       (n_4741));
  DFRQX1 \integer_file_reg[26][10] (.C (rc_gclk_205583), .D (n_62), .Q
       (n_5082));
  DFRQX1 \integer_file_reg[26][11] (.C (rc_gclk_205583), .D (n_77), .Q
       (n_5113));
  DFRQX1 \integer_file_reg[26][12] (.C (rc_gclk_205583), .D (n_38), .Q
       (n_5144));
  DFRQX1 \integer_file_reg[26][13] (.C (rc_gclk_205583), .D (n_54), .Q
       (n_5206));
  DFRQX1 \integer_file_reg[26][14] (.C (rc_gclk_205583), .D (n_37), .Q
       (n_5237));
  DFRQX1 \integer_file_reg[26][15] (.C (rc_gclk_205583), .D (n_53), .Q
       (n_5268));
  DFRQX1 \integer_file_reg[26][16] (.C (rc_gclk_205583), .D (n_65), .Q
       (n_5299));
  DFRQX1 \integer_file_reg[26][17] (.C (rc_gclk_205583), .D (n_75), .Q
       (n_5330));
  DFRQX1 \integer_file_reg[26][18] (.C (rc_gclk_205583), .D (n_43), .Q
       (n_5361));
  DFRQX1 \integer_file_reg[26][19] (.C (rc_gclk_205583), .D (n_51), .Q
       (n_5392));
  DFRQX1 \integer_file_reg[26][1] (.C (rc_gclk_205583), .D (n_15), .Q
       (n_4772));
  DFRQX1 \integer_file_reg[26][20] (.C (rc_gclk_205583), .D (n_60), .Q
       (n_5423));
  DFRQX1 \integer_file_reg[26][21] (.C (rc_gclk_205583), .D (n_59), .Q
       (n_5454));
  DFRQX1 \integer_file_reg[26][22] (.C (rc_gclk_205583), .D (n_56), .Q
       (n_5485));
  DFRQX1 \integer_file_reg[26][23] (.C (rc_gclk_205583), .D (n_71), .Q
       (n_4555));
  DFRQX1 \integer_file_reg[26][24] (.C (rc_gclk_205583), .D (n_64), .Q
       (n_4586));
  DFRQX1 \integer_file_reg[26][25] (.C (rc_gclk_205583), .D (n_36), .Q
       (n_4617));
  DFRQX1 \integer_file_reg[26][26] (.C (rc_gclk_205583), .D (n_31), .Q
       (n_4648));
  DFRQX1 \integer_file_reg[26][27] (.C (rc_gclk_205583), .D (n_69), .Q
       (n_4679));
  DFRQX1 \integer_file_reg[26][28] (.C (rc_gclk_205583), .D (n_41), .Q
       (n_4710));
  DFRQX1 \integer_file_reg[26][29] (.C (rc_gclk_205583), .D (n_42), .Q
       (n_4834));
  DFRQX1 \integer_file_reg[26][2] (.C (rc_gclk_205583), .D (n_16), .Q
       (n_4803));
  DFRQX1 \integer_file_reg[26][30] (.C (rc_gclk_205583), .D (n_48), .Q
       (n_5175));
  DFRQX1 \integer_file_reg[26][31] (.C (rc_gclk_205583), .D (n_68), .Q
       (n_5516));
  DFRQX1 \integer_file_reg[26][3] (.C (rc_gclk_205583), .D (n_25), .Q
       (n_4865));
  DFRQX1 \integer_file_reg[26][4] (.C (rc_gclk_205583), .D (n_22), .Q
       (n_4896));
  DFRQX1 \integer_file_reg[26][5] (.C (rc_gclk_205583), .D (n_30), .Q
       (n_4927));
  DFRQX1 \integer_file_reg[26][6] (.C (rc_gclk_205583), .D (n_20), .Q
       (n_4958));
  DFRQX1 \integer_file_reg[26][7] (.C (rc_gclk_205583), .D (n_33), .Q
       (n_4989));
  DFRQX1 \integer_file_reg[26][8] (.C (rc_gclk_205583), .D (n_67), .Q
       (n_5020));
  DFRQX1 \integer_file_reg[26][9] (.C (rc_gclk_205583), .D (n_47), .Q
       (n_5051));
  DFRQX1 \integer_file_reg[27][0] (.C (rc_gclk_205586), .D (n_26), .Q
       (n_4740));
  DFRQX1 \integer_file_reg[27][10] (.C (rc_gclk_205586), .D (n_78), .Q
       (n_5081));
  DFRQX1 \integer_file_reg[27][11] (.C (rc_gclk_205586), .D (n_66), .Q
       (n_5112));
  DFRQX1 \integer_file_reg[27][12] (.C (rc_gclk_205586), .D (n_28), .Q
       (n_5143));
  DFRQX1 \integer_file_reg[27][13] (.C (rc_gclk_205586), .D (n_44), .Q
       (n_5205));
  DFRQX1 \integer_file_reg[27][14] (.C (rc_gclk_205586), .D (n_37), .Q
       (n_5236));
  DFRQX1 \integer_file_reg[27][15] (.C (rc_gclk_205586), .D (n_53), .Q
       (n_5267));
  DFRQX1 \integer_file_reg[27][16] (.C (rc_gclk_205586), .D (n_65), .Q
       (n_5298));
  DFRQX1 \integer_file_reg[27][17] (.C (rc_gclk_205586), .D (n_75), .Q
       (n_5329));
  DFRQX1 \integer_file_reg[27][18] (.C (rc_gclk_205586), .D (n_43), .Q
       (n_5360));
  DFRQX1 \integer_file_reg[27][19] (.C (rc_gclk_205586), .D (n_39), .Q
       (n_5391));
  DFRQX1 \integer_file_reg[27][1] (.C (rc_gclk_205586), .D (n_15), .Q
       (n_4771));
  DFRQX1 \integer_file_reg[27][20] (.C (rc_gclk_205586), .D (n_74), .Q
       (n_5422));
  DFRQX1 \integer_file_reg[27][21] (.C (rc_gclk_205586), .D (n_73), .Q
       (n_5453));
  DFRQX1 \integer_file_reg[27][22] (.C (rc_gclk_205586), .D (n_56), .Q
       (n_5484));
  DFRQX1 \integer_file_reg[27][23] (.C (rc_gclk_205586), .D (n_55), .Q
       (n_4554));
  DFRQX1 \integer_file_reg[27][24] (.C (rc_gclk_205586), .D (n_70), .Q
       (n_4585));
  DFRQX1 \integer_file_reg[27][25] (.C (rc_gclk_205586), .D (n_27), .Q
       (n_4616));
  DFRQX1 \integer_file_reg[27][26] (.C (rc_gclk_205586), .D (n_31), .Q
       (n_4647));
  DFRQX1 \integer_file_reg[27][27] (.C (rc_gclk_205586), .D (n_69), .Q
       (n_4678));
  DFRQX1 \integer_file_reg[27][28] (.C (rc_gclk_205586), .D (n_41), .Q
       (n_4709));
  DFRQX1 \integer_file_reg[27][29] (.C (rc_gclk_205586), .D (n_42), .Q
       (n_4833));
  DFRQX1 \integer_file_reg[27][2] (.C (rc_gclk_205586), .D (n_17), .Q
       (n_4802));
  DFRQX1 \integer_file_reg[27][30] (.C (rc_gclk_205586), .D (n_48), .Q
       (n_5174));
  DFRQX1 \integer_file_reg[27][31] (.C (rc_gclk_205586), .D (n_63), .Q
       (n_5515));
  DFRQX1 \integer_file_reg[27][3] (.C (rc_gclk_205586), .D (n_25), .Q
       (n_4864));
  DFRQX1 \integer_file_reg[27][4] (.C (rc_gclk_205586), .D (n_22), .Q
       (n_4895));
  DFRQX1 \integer_file_reg[27][5] (.C (rc_gclk_205586), .D (n_30), .Q
       (n_4926));
  DFRQX1 \integer_file_reg[27][6] (.C (rc_gclk_205586), .D (n_23), .Q
       (n_4957));
  DFRQX1 \integer_file_reg[27][7] (.C (rc_gclk_205586), .D (n_33), .Q
       (n_4988));
  DFRQX1 \integer_file_reg[27][8] (.C (rc_gclk_205586), .D (n_57), .Q
       (n_5019));
  DFRQX1 \integer_file_reg[27][9] (.C (rc_gclk_205586), .D (n_40), .Q
       (n_5050));
  DFRQX1 \integer_file_reg[28][0] (.C (rc_gclk_205592), .D (n_26), .Q
       (n_4739));
  DFRQX1 \integer_file_reg[28][10] (.C (rc_gclk_205592), .D (n_78), .Q
       (n_5080));
  DFRQX1 \integer_file_reg[28][11] (.C (rc_gclk_205592), .D (n_66), .Q
       (n_5111));
  DFRQX1 \integer_file_reg[28][12] (.C (rc_gclk_205592), .D (n_38), .Q
       (n_5142));
  DFRQX1 \integer_file_reg[28][13] (.C (rc_gclk_205592), .D (n_44), .Q
       (n_5204));
  DFRQX1 \integer_file_reg[28][14] (.C (rc_gclk_205592), .D (n_37), .Q
       (n_5235));
  DFRQX1 \integer_file_reg[28][15] (.C (rc_gclk_205592), .D (n_53), .Q
       (n_5266));
  DFRQX1 \integer_file_reg[28][16] (.C (rc_gclk_205592), .D (n_65), .Q
       (n_5297));
  DFRQX1 \integer_file_reg[28][17] (.C (rc_gclk_205592), .D (n_75), .Q
       (n_5328));
  DFRQX1 \integer_file_reg[28][18] (.C (rc_gclk_205592), .D (n_52), .Q
       (n_5359));
  DFRQX1 \integer_file_reg[28][19] (.C (rc_gclk_205592), .D (n_51), .Q
       (n_5390));
  DFRQX1 \integer_file_reg[28][1] (.C (rc_gclk_205592), .D (n_15), .Q
       (n_4770));
  DFRQX1 \integer_file_reg[28][20] (.C (rc_gclk_205592), .D (n_74), .Q
       (n_5421));
  DFRQX1 \integer_file_reg[28][21] (.C (rc_gclk_205592), .D (n_73), .Q
       (n_5452));
  DFRQX1 \integer_file_reg[28][22] (.C (rc_gclk_205592), .D (n_72), .Q
       (n_5483));
  DFRQX1 \integer_file_reg[28][23] (.C (rc_gclk_205592), .D (n_71), .Q
       (n_4553));
  DFRQX1 \integer_file_reg[28][24] (.C (rc_gclk_205592), .D (n_64), .Q
       (n_4584));
  DFRQX1 \integer_file_reg[28][25] (.C (rc_gclk_205592), .D (n_27), .Q
       (n_4615));
  DFRQX1 \integer_file_reg[28][26] (.C (rc_gclk_205592), .D (n_35), .Q
       (n_4646));
  DFRQX1 \integer_file_reg[28][27] (.C (rc_gclk_205592), .D (n_69), .Q
       (n_4677));
  DFRQX1 \integer_file_reg[28][28] (.C (rc_gclk_205592), .D (n_50), .Q
       (n_4708));
  DFRQX1 \integer_file_reg[28][29] (.C (rc_gclk_205592), .D (n_49), .Q
       (n_4832));
  DFRQX1 \integer_file_reg[28][2] (.C (rc_gclk_205592), .D (n_17), .Q
       (n_4801));
  DFRQX1 \integer_file_reg[28][30] (.C (rc_gclk_205592), .D (n_48), .Q
       (n_5173));
  DFRQX1 \integer_file_reg[28][31] (.C (rc_gclk_205592), .D (n_68), .Q
       (n_5514));
  DFRQX1 \integer_file_reg[28][3] (.C (rc_gclk_205592), .D (n_19), .Q
       (n_4863));
  DFRQX1 \integer_file_reg[28][4] (.C (rc_gclk_205592), .D (n_22), .Q
       (n_4894));
  DFRQX1 \integer_file_reg[28][5] (.C (rc_gclk_205592), .D (n_34), .Q
       (n_4925));
  DFRQX1 \integer_file_reg[28][6] (.C (rc_gclk_205592), .D (n_20), .Q
       (n_4956));
  DFRQX1 \integer_file_reg[28][7] (.C (rc_gclk_205592), .D (n_29), .Q
       (n_4987));
  DFRQX1 \integer_file_reg[28][8] (.C (rc_gclk_205592), .D (n_57), .Q
       (n_5018));
  DFRQX1 \integer_file_reg[28][9] (.C (rc_gclk_205592), .D (n_47), .Q
       (n_5049));
  DFRQX1 \integer_file_reg[29][0] (.C (rc_gclk_205595), .D (n_26), .Q
       (n_4738));
  DFRQX1 \integer_file_reg[29][10] (.C (rc_gclk_205595), .D (n_78), .Q
       (n_5079));
  DFRQX1 \integer_file_reg[29][11] (.C (rc_gclk_205595), .D (n_66), .Q
       (n_5110));
  DFRQX1 \integer_file_reg[29][12] (.C (rc_gclk_205595), .D (n_38), .Q
       (n_5141));
  DFRQX1 \integer_file_reg[29][13] (.C (rc_gclk_205595), .D (n_44), .Q
       (n_5203));
  DFRQX1 \integer_file_reg[29][14] (.C (rc_gclk_205595), .D (n_37), .Q
       (n_5234));
  DFRQX1 \integer_file_reg[29][15] (.C (rc_gclk_205595), .D (n_53), .Q
       (n_5265));
  DFRQX1 \integer_file_reg[29][16] (.C (rc_gclk_205595), .D (n_76), .Q
       (n_5296));
  DFRQX1 \integer_file_reg[29][17] (.C (rc_gclk_205595), .D (n_61), .Q
       (n_5327));
  DFRQX1 \integer_file_reg[29][18] (.C (rc_gclk_205595), .D (n_43), .Q
       (n_5358));
  DFRQX1 \integer_file_reg[29][19] (.C (rc_gclk_205595), .D (n_51), .Q
       (n_5389));
  DFRQX1 \integer_file_reg[29][1] (.C (rc_gclk_205595), .D (n_18), .Q
       (n_4769));
  DFRQX1 \integer_file_reg[29][20] (.C (rc_gclk_205595), .D (n_60), .Q
       (n_5420));
  DFRQX1 \integer_file_reg[29][21] (.C (rc_gclk_205595), .D (n_73), .Q
       (n_5451));
  DFRQX1 \integer_file_reg[29][22] (.C (rc_gclk_205595), .D (n_72), .Q
       (n_5482));
  DFRQX1 \integer_file_reg[29][23] (.C (rc_gclk_205595), .D (n_71), .Q
       (n_4552));
  DFRQX1 \integer_file_reg[29][24] (.C (rc_gclk_205595), .D (n_70), .Q
       (n_4583));
  DFRQX1 \integer_file_reg[29][25] (.C (rc_gclk_205595), .D (n_36), .Q
       (n_4614));
  DFRQX1 \integer_file_reg[29][26] (.C (rc_gclk_205595), .D (n_35), .Q
       (n_4645));
  DFRQX1 \integer_file_reg[29][27] (.C (rc_gclk_205595), .D (n_58), .Q
       (n_4676));
  DFRQX1 \integer_file_reg[29][28] (.C (rc_gclk_205595), .D (n_50), .Q
       (n_4707));
  DFRQX1 \integer_file_reg[29][29] (.C (rc_gclk_205595), .D (n_49), .Q
       (n_4831));
  DFRQX1 \integer_file_reg[29][2] (.C (rc_gclk_205595), .D (n_16), .Q
       (n_4800));
  DFRQX1 \integer_file_reg[29][30] (.C (rc_gclk_205595), .D (n_45), .Q
       (n_5172));
  DFRQX1 \integer_file_reg[29][31] (.C (rc_gclk_205595), .D (n_68), .Q
       (n_5513));
  DFRQX1 \integer_file_reg[29][3] (.C (rc_gclk_205595), .D (n_25), .Q
       (n_4862));
  DFRQX1 \integer_file_reg[29][4] (.C (rc_gclk_205595), .D (n_24), .Q
       (n_4893));
  DFRQX1 \integer_file_reg[29][5] (.C (rc_gclk_205595), .D (n_34), .Q
       (n_4924));
  DFRQX1 \integer_file_reg[29][6] (.C (rc_gclk_205595), .D (n_23), .Q
       (n_4955));
  DFRQX1 \integer_file_reg[29][7] (.C (rc_gclk_205595), .D (n_33), .Q
       (n_4986));
  DFRQX1 \integer_file_reg[29][8] (.C (rc_gclk_205595), .D (n_67), .Q
       (n_5017));
  DFRQX1 \integer_file_reg[29][9] (.C (rc_gclk_205595), .D (n_47), .Q
       (n_5048));
  DFRQX1 \integer_file_reg[2][0] (.C (rc_gclk_205502), .D (n_21), .Q
       (n_4765));
  DFRQX1 \integer_file_reg[2][10] (.C (rc_gclk_205502), .D (n_78), .Q
       (n_5106));
  DFRQX1 \integer_file_reg[2][11] (.C (rc_gclk_205502), .D (n_66), .Q
       (n_5137));
  DFRQX1 \integer_file_reg[2][12] (.C (rc_gclk_205502), .D (n_38), .Q
       (n_5168));
  DFRQX1 \integer_file_reg[2][13] (.C (rc_gclk_205502), .D (n_54), .Q
       (n_5230));
  DFRQX1 \integer_file_reg[2][14] (.C (rc_gclk_205502), .D (n_32), .Q
       (n_5261));
  DFRQX1 \integer_file_reg[2][15] (.C (rc_gclk_205502), .D (n_53), .Q
       (n_5292));
  DFRQX1 \integer_file_reg[2][16] (.C (rc_gclk_205502), .D (n_65), .Q
       (n_5323));
  DFRQX1 \integer_file_reg[2][17] (.C (rc_gclk_205502), .D (n_61), .Q
       (n_5354));
  DFRQX1 \integer_file_reg[2][18] (.C (rc_gclk_205502), .D (n_43), .Q
       (n_5385));
  DFRQX1 \integer_file_reg[2][19] (.C (rc_gclk_205502), .D (n_51), .Q
       (n_5416));
  DFRQX1 \integer_file_reg[2][1] (.C (rc_gclk_205502), .D (n_15), .Q
       (n_4796));
  DFRQX1 \integer_file_reg[2][20] (.C (rc_gclk_205502), .D (n_60), .Q
       (n_5447));
  DFRQX1 \integer_file_reg[2][21] (.C (rc_gclk_205502), .D (n_73), .Q
       (n_5478));
  DFRQX1 \integer_file_reg[2][22] (.C (rc_gclk_205502), .D (n_72), .Q
       (n_5509));
  DFRQX1 \integer_file_reg[2][23] (.C (rc_gclk_205502), .D (n_71), .Q
       (n_4579));
  DFRQX1 \integer_file_reg[2][24] (.C (rc_gclk_205502), .D (n_64), .Q
       (n_4610));
  DFRQX1 \integer_file_reg[2][25] (.C (rc_gclk_205502), .D (n_27), .Q
       (n_4641));
  DFRQX1 \integer_file_reg[2][26] (.C (rc_gclk_205502), .D (n_31), .Q
       (n_4672));
  DFRQX1 \integer_file_reg[2][27] (.C (rc_gclk_205502), .D (n_69), .Q
       (n_4703));
  DFRQX1 \integer_file_reg[2][28] (.C (rc_gclk_205502), .D (n_50), .Q
       (n_4734));
  DFRQX1 \integer_file_reg[2][29] (.C (rc_gclk_205502), .D (n_49), .Q
       (n_4858));
  DFRQX1 \integer_file_reg[2][2] (.C (rc_gclk_205502), .D (n_17), .Q
       (n_4827));
  DFRQX1 \integer_file_reg[2][30] (.C (rc_gclk_205502), .D (n_48), .Q
       (n_5199));
  DFRQX1 \integer_file_reg[2][31] (.C (rc_gclk_205502), .D (n_63), .Q
       (n_5540));
  DFRQX1 \integer_file_reg[2][3] (.C (rc_gclk_205502), .D (n_25), .Q
       (n_4889));
  DFRQX1 \integer_file_reg[2][4] (.C (rc_gclk_205502), .D (n_22), .Q
       (n_4920));
  DFRQX1 \integer_file_reg[2][5] (.C (rc_gclk_205502), .D (n_34), .Q
       (n_4951));
  DFRQX1 \integer_file_reg[2][6] (.C (rc_gclk_205502), .D (n_23), .Q
       (n_4982));
  DFRQX1 \integer_file_reg[2][7] (.C (rc_gclk_205502), .D (n_33), .Q
       (n_5013));
  DFRQX1 \integer_file_reg[2][8] (.C (rc_gclk_205502), .D (n_67), .Q
       (n_5044));
  DFRQX1 \integer_file_reg[2][9] (.C (rc_gclk_205502), .D (n_40), .Q
       (n_5075));
  DFRQX1 \integer_file_reg[30][0] (.C (rc_gclk_205505), .D (n_21), .Q
       (n_4737));
  DFRQX1 \integer_file_reg[30][10] (.C (rc_gclk_205505), .D (n_78), .Q
       (n_5078));
  DFRQX1 \integer_file_reg[30][11] (.C (rc_gclk_205505), .D (n_66), .Q
       (n_5109));
  DFRQX1 \integer_file_reg[30][12] (.C (rc_gclk_205505), .D (n_38), .Q
       (n_5140));
  DFRQX1 \integer_file_reg[30][13] (.C (rc_gclk_205505), .D (n_44), .Q
       (n_5202));
  DFRQX1 \integer_file_reg[30][14] (.C (rc_gclk_205505), .D (n_37), .Q
       (n_5233));
  DFRQX1 \integer_file_reg[30][15] (.C (rc_gclk_205505), .D (n_53), .Q
       (n_5264));
  DFRQX1 \integer_file_reg[30][16] (.C (rc_gclk_205505), .D (n_76), .Q
       (n_5295));
  DFRQX1 \integer_file_reg[30][17] (.C (rc_gclk_205505), .D (n_61), .Q
       (n_5326));
  DFRQX1 \integer_file_reg[30][18] (.C (rc_gclk_205505), .D (n_43), .Q
       (n_5357));
  DFRQX1 \integer_file_reg[30][19] (.C (rc_gclk_205505), .D (n_39), .Q
       (n_5388));
  DFRQX1 \integer_file_reg[30][1] (.C (rc_gclk_205505), .D (n_18), .Q
       (n_4768));
  DFRQX1 \integer_file_reg[30][20] (.C (rc_gclk_205505), .D (n_60), .Q
       (n_5419));
  DFRQX1 \integer_file_reg[30][21] (.C (rc_gclk_205505), .D (n_59), .Q
       (n_5450));
  DFRQX1 \integer_file_reg[30][22] (.C (rc_gclk_205505), .D (n_56), .Q
       (n_5481));
  DFRQX1 \integer_file_reg[30][23] (.C (rc_gclk_205505), .D (n_55), .Q
       (n_4551));
  DFRQX1 \integer_file_reg[30][24] (.C (rc_gclk_205505), .D (n_64), .Q
       (n_4582));
  DFRQX1 \integer_file_reg[30][25] (.C (rc_gclk_205505), .D (n_36), .Q
       (n_4613));
  DFRQX1 \integer_file_reg[30][26] (.C (rc_gclk_205505), .D (n_35), .Q
       (n_4644));
  DFRQX1 \integer_file_reg[30][27] (.C (rc_gclk_205505), .D (n_69), .Q
       (n_4675));
  DFRQX1 \integer_file_reg[30][28] (.C (rc_gclk_205505), .D (n_50), .Q
       (n_4706));
  DFRQX1 \integer_file_reg[30][29] (.C (rc_gclk_205505), .D (n_49), .Q
       (n_4830));
  DFRQX1 \integer_file_reg[30][2] (.C (rc_gclk_205505), .D (n_17), .Q
       (n_4799));
  DFRQX1 \integer_file_reg[30][30] (.C (rc_gclk_205505), .D (n_45), .Q
       (n_5171));
  DFRQX1 \integer_file_reg[30][31] (.C (rc_gclk_205505), .D (n_63), .Q
       (n_5512));
  DFRQX1 \integer_file_reg[30][3] (.C (rc_gclk_205505), .D (n_25), .Q
       (n_4861));
  DFRQX1 \integer_file_reg[30][4] (.C (rc_gclk_205505), .D (n_22), .Q
       (n_4892));
  DFRQX1 \integer_file_reg[30][5] (.C (rc_gclk_205505), .D (n_34), .Q
       (n_4923));
  DFRQX1 \integer_file_reg[30][6] (.C (rc_gclk_205505), .D (n_23), .Q
       (n_4954));
  DFRQX1 \integer_file_reg[30][7] (.C (rc_gclk_205505), .D (n_33), .Q
       (n_4985));
  DFRQX1 \integer_file_reg[30][8] (.C (rc_gclk_205505), .D (n_67), .Q
       (n_5016));
  DFRQX1 \integer_file_reg[30][9] (.C (rc_gclk_205505), .D (n_47), .Q
       (n_5047));
  DFRQX1 \integer_file_reg[31][0] (.C (rc_gclk_205511), .D (n_26), .Q
       (n_4736));
  DFRQX1 \integer_file_reg[31][10] (.C (rc_gclk_205511), .D (n_78), .Q
       (n_5077));
  DFRQX1 \integer_file_reg[31][11] (.C (rc_gclk_205511), .D (n_66), .Q
       (n_5108));
  DFRQX1 \integer_file_reg[31][12] (.C (rc_gclk_205511), .D (n_28), .Q
       (n_5139));
  DFRQX1 \integer_file_reg[31][13] (.C (rc_gclk_205511), .D (n_44), .Q
       (n_5201));
  DFRQX1 \integer_file_reg[31][14] (.C (rc_gclk_205511), .D (n_37), .Q
       (n_5232));
  DFRQX1 \integer_file_reg[31][15] (.C (rc_gclk_205511), .D (n_53), .Q
       (n_5263));
  DFRQX1 \integer_file_reg[31][16] (.C (rc_gclk_205511), .D (n_65), .Q
       (n_5294));
  DFRQX1 \integer_file_reg[31][17] (.C (rc_gclk_205511), .D (n_75), .Q
       (n_5325));
  DFRQX1 \integer_file_reg[31][18] (.C (rc_gclk_205511), .D (n_43), .Q
       (n_5356));
  DFRQX1 \integer_file_reg[31][19] (.C (rc_gclk_205511), .D (n_51), .Q
       (n_5387));
  DFRQX1 \integer_file_reg[31][1] (.C (rc_gclk_205511), .D (n_18), .Q
       (n_4767));
  DFRQX1 \integer_file_reg[31][20] (.C (rc_gclk_205511), .D (n_74), .Q
       (n_5418));
  DFRQX1 \integer_file_reg[31][21] (.C (rc_gclk_205511), .D (n_73), .Q
       (n_5449));
  DFRQX1 \integer_file_reg[31][22] (.C (rc_gclk_205511), .D (n_56), .Q
       (n_5480));
  DFRQX1 \integer_file_reg[31][23] (.C (rc_gclk_205511), .D (n_71), .Q
       (n_4550));
  DFRQX1 \integer_file_reg[31][24] (.C (rc_gclk_205511), .D (n_64), .Q
       (n_4581));
  DFRQX1 \integer_file_reg[31][25] (.C (rc_gclk_205511), .D (n_27), .Q
       (n_4612));
  DFRQX1 \integer_file_reg[31][26] (.C (rc_gclk_205511), .D (n_31), .Q
       (n_4643));
  DFRQX1 \integer_file_reg[31][27] (.C (rc_gclk_205511), .D (n_69), .Q
       (n_4674));
  DFRQX1 \integer_file_reg[31][28] (.C (rc_gclk_205511), .D (n_41), .Q
       (n_4705));
  DFRQX1 \integer_file_reg[31][29] (.C (rc_gclk_205511), .D (n_49), .Q
       (n_4829));
  DFRQX1 \integer_file_reg[31][2] (.C (rc_gclk_205511), .D (n_17), .Q
       (n_4798));
  DFRQX1 \integer_file_reg[31][30] (.C (rc_gclk_205511), .D (n_45), .Q
       (n_5170));
  DFRQX1 \integer_file_reg[31][31] (.C (rc_gclk_205511), .D (n_63), .Q
       (n_5511));
  DFRQX1 \integer_file_reg[31][3] (.C (rc_gclk_205511), .D (n_25), .Q
       (n_4860));
  DFRQX1 \integer_file_reg[31][4] (.C (rc_gclk_205511), .D (n_24), .Q
       (n_4891));
  DFRQX1 \integer_file_reg[31][5] (.C (rc_gclk_205511), .D (n_34), .Q
       (n_4922));
  DFRQX1 \integer_file_reg[31][6] (.C (rc_gclk_205511), .D (n_23), .Q
       (n_4953));
  DFRQX1 \integer_file_reg[31][7] (.C (rc_gclk_205511), .D (n_29), .Q
       (n_4984));
  DFRQX1 \integer_file_reg[31][8] (.C (rc_gclk_205511), .D (n_57), .Q
       (n_5015));
  DFRQX1 \integer_file_reg[31][9] (.C (rc_gclk_205511), .D (n_40), .Q
       (n_5046));
  DFRQX1 \integer_file_reg[3][0] (.C (rc_gclk_205514), .D (n_21), .Q
       (n_4764));
  DFRQX1 \integer_file_reg[3][10] (.C (rc_gclk_205514), .D (n_62), .Q
       (n_5105));
  DFRQX1 \integer_file_reg[3][11] (.C (rc_gclk_205514), .D (n_77), .Q
       (n_5136));
  DFRQX1 \integer_file_reg[3][12] (.C (rc_gclk_205514), .D (n_28), .Q
       (n_5167));
  DFRQX1 \integer_file_reg[3][13] (.C (rc_gclk_205514), .D (n_54), .Q
       (n_5229));
  DFRQX1 \integer_file_reg[3][14] (.C (rc_gclk_205514), .D (n_37), .Q
       (n_5260));
  DFRQX1 \integer_file_reg[3][15] (.C (rc_gclk_205514), .D (n_53), .Q
       (n_5291));
  DFRQX1 \integer_file_reg[3][16] (.C (rc_gclk_205514), .D (n_65), .Q
       (n_5322));
  DFRQX1 \integer_file_reg[3][17] (.C (rc_gclk_205514), .D (n_75), .Q
       (n_5353));
  DFRQX1 \integer_file_reg[3][18] (.C (rc_gclk_205514), .D (n_52), .Q
       (n_5384));
  DFRQX1 \integer_file_reg[3][19] (.C (rc_gclk_205514), .D (n_51), .Q
       (n_5415));
  DFRQX1 \integer_file_reg[3][1] (.C (rc_gclk_205514), .D (n_15), .Q
       (n_4795));
  DFRQX1 \integer_file_reg[3][20] (.C (rc_gclk_205514), .D (n_60), .Q
       (n_5446));
  DFRQX1 \integer_file_reg[3][21] (.C (rc_gclk_205514), .D (n_73), .Q
       (n_5477));
  DFRQX1 \integer_file_reg[3][22] (.C (rc_gclk_205514), .D (n_56), .Q
       (n_5508));
  DFRQX1 \integer_file_reg[3][23] (.C (rc_gclk_205514), .D (n_71), .Q
       (n_4578));
  DFRQX1 \integer_file_reg[3][24] (.C (rc_gclk_205514), .D (n_64), .Q
       (n_4609));
  DFRQX1 \integer_file_reg[3][25] (.C (rc_gclk_205514), .D (n_36), .Q
       (n_4640));
  DFRQX1 \integer_file_reg[3][26] (.C (rc_gclk_205514), .D (n_31), .Q
       (n_4671));
  DFRQX1 \integer_file_reg[3][27] (.C (rc_gclk_205514), .D (n_69), .Q
       (n_4702));
  DFRQX1 \integer_file_reg[3][28] (.C (rc_gclk_205514), .D (n_50), .Q
       (n_4733));
  DFRQX1 \integer_file_reg[3][29] (.C (rc_gclk_205514), .D (n_49), .Q
       (n_4857));
  DFRQX1 \integer_file_reg[3][2] (.C (rc_gclk_205514), .D (n_17), .Q
       (n_4826));
  DFRQX1 \integer_file_reg[3][30] (.C (rc_gclk_205514), .D (n_45), .Q
       (n_5198));
  DFRQX1 \integer_file_reg[3][31] (.C (rc_gclk_205514), .D (n_63), .Q
       (n_5539));
  DFRQX1 \integer_file_reg[3][3] (.C (rc_gclk_205514), .D (n_25), .Q
       (n_4888));
  DFRQX1 \integer_file_reg[3][4] (.C (rc_gclk_205514), .D (n_24), .Q
       (n_4919));
  DFRQX1 \integer_file_reg[3][5] (.C (rc_gclk_205514), .D (n_34), .Q
       (n_4950));
  DFRQX1 \integer_file_reg[3][6] (.C (rc_gclk_205514), .D (n_23), .Q
       (n_4981));
  DFRQX1 \integer_file_reg[3][7] (.C (rc_gclk_205514), .D (n_33), .Q
       (n_5012));
  DFRQX1 \integer_file_reg[3][8] (.C (rc_gclk_205514), .D (n_67), .Q
       (n_5043));
  DFRQX1 \integer_file_reg[3][9] (.C (rc_gclk_205514), .D (n_47), .Q
       (n_5074));
  DFRQX1 \integer_file_reg[4][0] (.C (rc_gclk_205520), .D (n_26), .Q
       (n_4763));
  DFRQX1 \integer_file_reg[4][10] (.C (rc_gclk_205520), .D (n_62), .Q
       (n_5104));
  DFRQX1 \integer_file_reg[4][11] (.C (rc_gclk_205520), .D (n_66), .Q
       (n_5135));
  DFRQX1 \integer_file_reg[4][12] (.C (rc_gclk_205520), .D (n_28), .Q
       (n_5166));
  DFRQX1 \integer_file_reg[4][13] (.C (rc_gclk_205520), .D (n_44), .Q
       (n_5228));
  DFRQX1 \integer_file_reg[4][14] (.C (rc_gclk_205520), .D (n_37), .Q
       (n_5259));
  DFRQX1 \integer_file_reg[4][15] (.C (rc_gclk_205520), .D (n_53), .Q
       (n_5290));
  DFRQX1 \integer_file_reg[4][16] (.C (rc_gclk_205520), .D (n_65), .Q
       (n_5321));
  DFRQX1 \integer_file_reg[4][17] (.C (rc_gclk_205520), .D (n_61), .Q
       (n_5352));
  DFRQX1 \integer_file_reg[4][18] (.C (rc_gclk_205520), .D (n_43), .Q
       (n_5383));
  DFRQX1 \integer_file_reg[4][19] (.C (rc_gclk_205520), .D (n_51), .Q
       (n_5414));
  DFRQX1 \integer_file_reg[4][1] (.C (rc_gclk_205520), .D (n_15), .Q
       (n_4794));
  DFRQX1 \integer_file_reg[4][20] (.C (rc_gclk_205520), .D (n_74), .Q
       (n_5445));
  DFRQX1 \integer_file_reg[4][21] (.C (rc_gclk_205520), .D (n_59), .Q
       (n_5476));
  DFRQX1 \integer_file_reg[4][22] (.C (rc_gclk_205520), .D (n_72), .Q
       (n_5507));
  DFRQX1 \integer_file_reg[4][23] (.C (rc_gclk_205520), .D (n_71), .Q
       (n_4577));
  DFRQX1 \integer_file_reg[4][24] (.C (rc_gclk_205520), .D (n_64), .Q
       (n_4608));
  DFRQX1 \integer_file_reg[4][25] (.C (rc_gclk_205520), .D (n_36), .Q
       (n_4639));
  DFRQX1 \integer_file_reg[4][26] (.C (rc_gclk_205520), .D (n_31), .Q
       (n_4670));
  DFRQX1 \integer_file_reg[4][27] (.C (rc_gclk_205520), .D (n_58), .Q
       (n_4701));
  DFRQX1 \integer_file_reg[4][28] (.C (rc_gclk_205520), .D (n_50), .Q
       (n_4732));
  DFRQX1 \integer_file_reg[4][29] (.C (rc_gclk_205520), .D (n_49), .Q
       (n_4856));
  DFRQX1 \integer_file_reg[4][2] (.C (rc_gclk_205520), .D (n_17), .Q
       (n_4825));
  DFRQX1 \integer_file_reg[4][30] (.C (rc_gclk_205520), .D (n_48), .Q
       (n_5197));
  DFRQX1 \integer_file_reg[4][31] (.C (rc_gclk_205520), .D (n_63), .Q
       (n_5538));
  DFRQX1 \integer_file_reg[4][3] (.C (rc_gclk_205520), .D (n_25), .Q
       (n_4887));
  DFRQX1 \integer_file_reg[4][4] (.C (rc_gclk_205520), .D (n_24), .Q
       (n_4918));
  DFRQX1 \integer_file_reg[4][5] (.C (rc_gclk_205520), .D (n_34), .Q
       (n_4949));
  DFRQX1 \integer_file_reg[4][6] (.C (rc_gclk_205520), .D (n_23), .Q
       (n_4980));
  DFRQX1 \integer_file_reg[4][7] (.C (rc_gclk_205520), .D (n_33), .Q
       (n_5011));
  DFRQX1 \integer_file_reg[4][8] (.C (rc_gclk_205520), .D (n_67), .Q
       (n_5042));
  DFRQX1 \integer_file_reg[4][9] (.C (rc_gclk_205520), .D (n_47), .Q
       (n_5073));
  DFRQX1 \integer_file_reg[5][0] (.C (rc_gclk_205523), .D (n_26), .Q
       (n_4762));
  DFRQX1 \integer_file_reg[5][10] (.C (rc_gclk_205523), .D (n_78), .Q
       (n_5103));
  DFRQX1 \integer_file_reg[5][11] (.C (rc_gclk_205523), .D (n_66), .Q
       (n_5134));
  DFRQX1 \integer_file_reg[5][12] (.C (rc_gclk_205523), .D (n_38), .Q
       (n_5165));
  DFRQX1 \integer_file_reg[5][13] (.C (rc_gclk_205523), .D (n_54), .Q
       (n_5227));
  DFRQX1 \integer_file_reg[5][14] (.C (rc_gclk_205523), .D (n_37), .Q
       (n_5258));
  DFRQX1 \integer_file_reg[5][15] (.C (rc_gclk_205523), .D (n_53), .Q
       (n_5289));
  DFRQX1 \integer_file_reg[5][16] (.C (rc_gclk_205523), .D (n_65), .Q
       (n_5320));
  DFRQX1 \integer_file_reg[5][17] (.C (rc_gclk_205523), .D (n_61), .Q
       (n_5351));
  DFRQX1 \integer_file_reg[5][18] (.C (rc_gclk_205523), .D (n_52), .Q
       (n_5382));
  DFRQX1 \integer_file_reg[5][19] (.C (rc_gclk_205523), .D (n_51), .Q
       (n_5413));
  DFRQX1 \integer_file_reg[5][1] (.C (rc_gclk_205523), .D (n_15), .Q
       (n_4793));
  DFRQX1 \integer_file_reg[5][20] (.C (rc_gclk_205523), .D (n_60), .Q
       (n_5444));
  DFRQX1 \integer_file_reg[5][21] (.C (rc_gclk_205523), .D (n_59), .Q
       (n_5475));
  DFRQX1 \integer_file_reg[5][22] (.C (rc_gclk_205523), .D (n_72), .Q
       (n_5506));
  DFRQX1 \integer_file_reg[5][23] (.C (rc_gclk_205523), .D (n_55), .Q
       (n_4576));
  DFRQX1 \integer_file_reg[5][24] (.C (rc_gclk_205523), .D (n_64), .Q
       (n_4607));
  DFRQX1 \integer_file_reg[5][25] (.C (rc_gclk_205523), .D (n_36), .Q
       (n_4638));
  DFRQX1 \integer_file_reg[5][26] (.C (rc_gclk_205523), .D (n_31), .Q
       (n_4669));
  DFRQX1 \integer_file_reg[5][27] (.C (rc_gclk_205523), .D (n_69), .Q
       (n_4700));
  DFRQX1 \integer_file_reg[5][28] (.C (rc_gclk_205523), .D (n_50), .Q
       (n_4731));
  DFRQX1 \integer_file_reg[5][29] (.C (rc_gclk_205523), .D (n_42), .Q
       (n_4855));
  DFRQX1 \integer_file_reg[5][2] (.C (rc_gclk_205523), .D (n_16), .Q
       (n_4824));
  DFRQX1 \integer_file_reg[5][30] (.C (rc_gclk_205523), .D (n_45), .Q
       (n_5196));
  DFRQX1 \integer_file_reg[5][31] (.C (rc_gclk_205523), .D (n_63), .Q
       (n_5537));
  DFRQX1 \integer_file_reg[5][3] (.C (rc_gclk_205523), .D (n_25), .Q
       (n_4886));
  DFRQX1 \integer_file_reg[5][4] (.C (rc_gclk_205523), .D (n_22), .Q
       (n_4917));
  DFRQX1 \integer_file_reg[5][5] (.C (rc_gclk_205523), .D (n_34), .Q
       (n_4948));
  DFRQX1 \integer_file_reg[5][6] (.C (rc_gclk_205523), .D (n_23), .Q
       (n_4979));
  DFRQX1 \integer_file_reg[5][7] (.C (rc_gclk_205523), .D (n_33), .Q
       (n_5010));
  DFRQX1 \integer_file_reg[5][8] (.C (rc_gclk_205523), .D (n_67), .Q
       (n_5041));
  DFRQX1 \integer_file_reg[5][9] (.C (rc_gclk_205523), .D (n_47), .Q
       (n_5072));
  DFRQX1 \integer_file_reg[6][0] (.C (rc_gclk_205529), .D (n_26), .Q
       (n_4761));
  DFRQX1 \integer_file_reg[6][10] (.C (rc_gclk_205529), .D (n_78), .Q
       (n_5102));
  DFRQX1 \integer_file_reg[6][11] (.C (rc_gclk_205529), .D (n_77), .Q
       (n_5133));
  DFRQX1 \integer_file_reg[6][12] (.C (rc_gclk_205529), .D (n_38), .Q
       (n_5164));
  DFRQX1 \integer_file_reg[6][13] (.C (rc_gclk_205529), .D (n_54), .Q
       (n_5226));
  DFRQX1 \integer_file_reg[6][14] (.C (rc_gclk_205529), .D (n_37), .Q
       (n_5257));
  DFRQX1 \integer_file_reg[6][15] (.C (rc_gclk_205529), .D (n_46), .Q
       (n_5288));
  DFRQX1 \integer_file_reg[6][16] (.C (rc_gclk_205529), .D (n_65), .Q
       (n_5319));
  DFRQX1 \integer_file_reg[6][17] (.C (rc_gclk_205529), .D (n_75), .Q
       (n_5350));
  DFRQX1 \integer_file_reg[6][18] (.C (rc_gclk_205529), .D (n_52), .Q
       (n_5381));
  DFRQX1 \integer_file_reg[6][19] (.C (rc_gclk_205529), .D (n_51), .Q
       (n_5412));
  DFRQX1 \integer_file_reg[6][1] (.C (rc_gclk_205529), .D (n_18), .Q
       (n_4792));
  DFRQX1 \integer_file_reg[6][20] (.C (rc_gclk_205529), .D (n_74), .Q
       (n_5443));
  DFRQX1 \integer_file_reg[6][21] (.C (rc_gclk_205529), .D (n_73), .Q
       (n_5474));
  DFRQX1 \integer_file_reg[6][22] (.C (rc_gclk_205529), .D (n_56), .Q
       (n_5505));
  DFRQX1 \integer_file_reg[6][23] (.C (rc_gclk_205529), .D (n_55), .Q
       (n_4575));
  DFRQX1 \integer_file_reg[6][24] (.C (rc_gclk_205529), .D (n_64), .Q
       (n_4606));
  DFRQX1 \integer_file_reg[6][25] (.C (rc_gclk_205529), .D (n_36), .Q
       (n_4637));
  DFRQX1 \integer_file_reg[6][26] (.C (rc_gclk_205529), .D (n_31), .Q
       (n_4668));
  DFRQX1 \integer_file_reg[6][27] (.C (rc_gclk_205529), .D (n_69), .Q
       (n_4699));
  DFRQX1 \integer_file_reg[6][28] (.C (rc_gclk_205529), .D (n_41), .Q
       (n_4730));
  DFRQX1 \integer_file_reg[6][29] (.C (rc_gclk_205529), .D (n_42), .Q
       (n_4854));
  DFRQX1 \integer_file_reg[6][2] (.C (rc_gclk_205529), .D (n_17), .Q
       (n_4823));
  DFRQX1 \integer_file_reg[6][30] (.C (rc_gclk_205529), .D (n_45), .Q
       (n_5195));
  DFRQX1 \integer_file_reg[6][31] (.C (rc_gclk_205529), .D (n_63), .Q
       (n_5536));
  DFRQX1 \integer_file_reg[6][3] (.C (rc_gclk_205529), .D (n_25), .Q
       (n_4885));
  DFRQX1 \integer_file_reg[6][4] (.C (rc_gclk_205529), .D (n_22), .Q
       (n_4916));
  DFRQX1 \integer_file_reg[6][5] (.C (rc_gclk_205529), .D (n_34), .Q
       (n_4947));
  DFRQX1 \integer_file_reg[6][6] (.C (rc_gclk_205529), .D (n_23), .Q
       (n_4978));
  DFRQX1 \integer_file_reg[6][7] (.C (rc_gclk_205529), .D (n_33), .Q
       (n_5009));
  DFRQX1 \integer_file_reg[6][8] (.C (rc_gclk_205529), .D (n_57), .Q
       (n_5040));
  DFRQX1 \integer_file_reg[6][9] (.C (rc_gclk_205529), .D (n_47), .Q
       (n_5071));
  DFRQX1 \integer_file_reg[7][0] (.C (rc_gclk_205532), .D (n_26), .Q
       (n_4760));
  DFRQX1 \integer_file_reg[7][10] (.C (rc_gclk_205532), .D (n_78), .Q
       (n_5101));
  DFRQX1 \integer_file_reg[7][11] (.C (rc_gclk_205532), .D (n_66), .Q
       (n_5132));
  DFRQX1 \integer_file_reg[7][12] (.C (rc_gclk_205532), .D (n_38), .Q
       (n_5163));
  DFRQX1 \integer_file_reg[7][13] (.C (rc_gclk_205532), .D (n_44), .Q
       (n_5225));
  DFRQX1 \integer_file_reg[7][14] (.C (rc_gclk_205532), .D (n_37), .Q
       (n_5256));
  DFRQX1 \integer_file_reg[7][15] (.C (rc_gclk_205532), .D (n_53), .Q
       (n_5287));
  DFRQX1 \integer_file_reg[7][16] (.C (rc_gclk_205532), .D (n_76), .Q
       (n_5318));
  DFRQX1 \integer_file_reg[7][17] (.C (rc_gclk_205532), .D (n_61), .Q
       (n_5349));
  DFRQX1 \integer_file_reg[7][18] (.C (rc_gclk_205532), .D (n_52), .Q
       (n_5380));
  DFRQX1 \integer_file_reg[7][19] (.C (rc_gclk_205532), .D (n_39), .Q
       (n_5411));
  DFRQX1 \integer_file_reg[7][1] (.C (rc_gclk_205532), .D (n_15), .Q
       (n_4791));
  DFRQX1 \integer_file_reg[7][20] (.C (rc_gclk_205532), .D (n_74), .Q
       (n_5442));
  DFRQX1 \integer_file_reg[7][21] (.C (rc_gclk_205532), .D (n_59), .Q
       (n_5473));
  DFRQX1 \integer_file_reg[7][22] (.C (rc_gclk_205532), .D (n_56), .Q
       (n_5504));
  DFRQX1 \integer_file_reg[7][23] (.C (rc_gclk_205532), .D (n_55), .Q
       (n_4574));
  DFRQX1 \integer_file_reg[7][24] (.C (rc_gclk_205532), .D (n_64), .Q
       (n_4605));
  DFRQX1 \integer_file_reg[7][25] (.C (rc_gclk_205532), .D (n_27), .Q
       (n_4636));
  DFRQX1 \integer_file_reg[7][26] (.C (rc_gclk_205532), .D (n_35), .Q
       (n_4667));
  DFRQX1 \integer_file_reg[7][27] (.C (rc_gclk_205532), .D (n_69), .Q
       (n_4698));
  DFRQX1 \integer_file_reg[7][28] (.C (rc_gclk_205532), .D (n_50), .Q
       (n_4729));
  DFRQX1 \integer_file_reg[7][29] (.C (rc_gclk_205532), .D (n_42), .Q
       (n_4853));
  DFRQX1 \integer_file_reg[7][2] (.C (rc_gclk_205532), .D (n_17), .Q
       (n_4822));
  DFRQX1 \integer_file_reg[7][30] (.C (rc_gclk_205532), .D (n_45), .Q
       (n_5194));
  DFRQX1 \integer_file_reg[7][31] (.C (rc_gclk_205532), .D (n_63), .Q
       (n_5535));
  DFRQX1 \integer_file_reg[7][3] (.C (rc_gclk_205532), .D (n_25), .Q
       (n_4884));
  DFRQX1 \integer_file_reg[7][4] (.C (rc_gclk_205532), .D (n_22), .Q
       (n_4915));
  DFRQX1 \integer_file_reg[7][5] (.C (rc_gclk_205532), .D (n_34), .Q
       (n_4946));
  DFRQX1 \integer_file_reg[7][6] (.C (rc_gclk_205532), .D (n_23), .Q
       (n_4977));
  DFRQX1 \integer_file_reg[7][7] (.C (rc_gclk_205532), .D (n_33), .Q
       (n_5008));
  DFRQX1 \integer_file_reg[7][8] (.C (rc_gclk_205532), .D (n_67), .Q
       (n_5039));
  DFRQX1 \integer_file_reg[7][9] (.C (rc_gclk_205532), .D (n_47), .Q
       (n_5070));
  DFRQX1 \integer_file_reg[8][0] (.C (rc_gclk_205541), .D (n_26), .Q
       (n_4759));
  DFRQX1 \integer_file_reg[8][10] (.C (rc_gclk_205541), .D (n_62), .Q
       (n_5100));
  DFRQX1 \integer_file_reg[8][11] (.C (rc_gclk_205541), .D (n_66), .Q
       (n_5131));
  DFRQX1 \integer_file_reg[8][12] (.C (rc_gclk_205541), .D (n_38), .Q
       (n_5162));
  DFRQX1 \integer_file_reg[8][13] (.C (rc_gclk_205541), .D (n_44), .Q
       (n_5224));
  DFRQX1 \integer_file_reg[8][14] (.C (rc_gclk_205541), .D (n_37), .Q
       (n_5255));
  DFRQX1 \integer_file_reg[8][15] (.C (rc_gclk_205541), .D (n_46), .Q
       (n_5286));
  DFRQX1 \integer_file_reg[8][16] (.C (rc_gclk_205541), .D (n_76), .Q
       (n_5317));
  DFRQX1 \integer_file_reg[8][17] (.C (rc_gclk_205541), .D (n_75), .Q
       (n_5348));
  DFRQX1 \integer_file_reg[8][18] (.C (rc_gclk_205541), .D (n_43), .Q
       (n_5379));
  DFRQX1 \integer_file_reg[8][19] (.C (rc_gclk_205541), .D (n_51), .Q
       (n_5410));
  DFRQX1 \integer_file_reg[8][1] (.C (rc_gclk_205541), .D (n_18), .Q
       (n_4790));
  DFRQX1 \integer_file_reg[8][20] (.C (rc_gclk_205541), .D (n_60), .Q
       (n_5441));
  DFRQX1 \integer_file_reg[8][21] (.C (rc_gclk_205541), .D (n_73), .Q
       (n_5472));
  DFRQX1 \integer_file_reg[8][22] (.C (rc_gclk_205541), .D (n_72), .Q
       (n_5503));
  DFRQX1 \integer_file_reg[8][23] (.C (rc_gclk_205541), .D (n_55), .Q
       (n_4573));
  DFRQX1 \integer_file_reg[8][24] (.C (rc_gclk_205541), .D (n_64), .Q
       (n_4604));
  DFRQX1 \integer_file_reg[8][25] (.C (rc_gclk_205541), .D (n_27), .Q
       (n_4635));
  DFRQX1 \integer_file_reg[8][26] (.C (rc_gclk_205541), .D (n_31), .Q
       (n_4666));
  DFRQX1 \integer_file_reg[8][27] (.C (rc_gclk_205541), .D (n_69), .Q
       (n_4697));
  DFRQX1 \integer_file_reg[8][28] (.C (rc_gclk_205541), .D (n_41), .Q
       (n_4728));
  DFRQX1 \integer_file_reg[8][29] (.C (rc_gclk_205541), .D (n_49), .Q
       (n_4852));
  DFRQX1 \integer_file_reg[8][2] (.C (rc_gclk_205541), .D (n_16), .Q
       (n_4821));
  DFRQX1 \integer_file_reg[8][30] (.C (rc_gclk_205541), .D (n_48), .Q
       (n_5193));
  DFRQX1 \integer_file_reg[8][31] (.C (rc_gclk_205541), .D (n_68), .Q
       (n_5534));
  DFRQX1 \integer_file_reg[8][3] (.C (rc_gclk_205541), .D (n_19), .Q
       (n_4883));
  DFRQX1 \integer_file_reg[8][4] (.C (rc_gclk_205541), .D (n_22), .Q
       (n_4914));
  DFRQX1 \integer_file_reg[8][5] (.C (rc_gclk_205541), .D (n_34), .Q
       (n_4945));
  DFRQX1 \integer_file_reg[8][6] (.C (rc_gclk_205541), .D (n_23), .Q
       (n_4976));
  DFRQX1 \integer_file_reg[8][7] (.C (rc_gclk_205541), .D (n_29), .Q
       (n_5007));
  DFRQX1 \integer_file_reg[8][8] (.C (rc_gclk_205541), .D (n_67), .Q
       (n_5038));
  DFRQX1 \integer_file_reg[8][9] (.C (rc_gclk_205541), .D (n_47), .Q
       (n_5069));
  DFRQX1 \integer_file_reg[9][0] (.C (rc_gclk_205544), .D (n_26), .Q
       (n_4758));
  DFRQX1 \integer_file_reg[9][10] (.C (rc_gclk_205544), .D (n_62), .Q
       (n_5099));
  DFRQX1 \integer_file_reg[9][11] (.C (rc_gclk_205544), .D (n_77), .Q
       (n_5130));
  DFRQX1 \integer_file_reg[9][12] (.C (rc_gclk_205544), .D (n_38), .Q
       (n_5161));
  DFRQX1 \integer_file_reg[9][13] (.C (rc_gclk_205544), .D (n_44), .Q
       (n_5223));
  DFRQX1 \integer_file_reg[9][14] (.C (rc_gclk_205544), .D (n_37), .Q
       (n_5254));
  DFRQX1 \integer_file_reg[9][15] (.C (rc_gclk_205544), .D (n_53), .Q
       (n_5285));
  DFRQX1 \integer_file_reg[9][16] (.C (rc_gclk_205544), .D (n_65), .Q
       (n_5316));
  DFRQX1 \integer_file_reg[9][17] (.C (rc_gclk_205544), .D (n_61), .Q
       (n_5347));
  DFRQX1 \integer_file_reg[9][18] (.C (rc_gclk_205544), .D (n_52), .Q
       (n_5378));
  DFRQX1 \integer_file_reg[9][19] (.C (rc_gclk_205544), .D (n_51), .Q
       (n_5409));
  DFRQX1 \integer_file_reg[9][1] (.C (rc_gclk_205544), .D (n_15), .Q
       (n_4789));
  DFRQX1 \integer_file_reg[9][20] (.C (rc_gclk_205544), .D (n_60), .Q
       (n_5440));
  DFRQX1 \integer_file_reg[9][21] (.C (rc_gclk_205544), .D (n_73), .Q
       (n_5471));
  DFRQX1 \integer_file_reg[9][22] (.C (rc_gclk_205544), .D (n_72), .Q
       (n_5502));
  DFRQX1 \integer_file_reg[9][23] (.C (rc_gclk_205544), .D (n_71), .Q
       (n_4572));
  DFRQX1 \integer_file_reg[9][24] (.C (rc_gclk_205544), .D (n_64), .Q
       (n_4603));
  DFRQX1 \integer_file_reg[9][25] (.C (rc_gclk_205544), .D (n_36), .Q
       (n_4634));
  DFRQX1 \integer_file_reg[9][26] (.C (rc_gclk_205544), .D (n_31), .Q
       (n_4665));
  DFRQX1 \integer_file_reg[9][27] (.C (rc_gclk_205544), .D (n_69), .Q
       (n_4696));
  DFRQX1 \integer_file_reg[9][28] (.C (rc_gclk_205544), .D (n_50), .Q
       (n_4727));
  DFRQX1 \integer_file_reg[9][29] (.C (rc_gclk_205544), .D (n_42), .Q
       (n_4851));
  DFRQX1 \integer_file_reg[9][2] (.C (rc_gclk_205544), .D (n_17), .Q
       (n_4820));
  DFRQX1 \integer_file_reg[9][30] (.C (rc_gclk_205544), .D (n_48), .Q
       (n_5192));
  DFRQX1 \integer_file_reg[9][31] (.C (rc_gclk_205544), .D (n_68), .Q
       (n_5533));
  DFRQX1 \integer_file_reg[9][3] (.C (rc_gclk_205544), .D (n_25), .Q
       (n_4882));
  DFRQX1 \integer_file_reg[9][4] (.C (rc_gclk_205544), .D (n_24), .Q
       (n_4913));
  DFRQX1 \integer_file_reg[9][5] (.C (rc_gclk_205544), .D (n_34), .Q
       (n_4944));
  DFRQX1 \integer_file_reg[9][6] (.C (rc_gclk_205544), .D (n_23), .Q
       (n_4975));
  DFRQX1 \integer_file_reg[9][7] (.C (rc_gclk_205544), .D (n_33), .Q
       (n_5006));
  DFRQX1 \integer_file_reg[9][8] (.C (rc_gclk_205544), .D (n_57), .Q
       (n_5037));
  DFRQX1 \integer_file_reg[9][9] (.C (rc_gclk_205544), .D (n_40), .Q
       (n_5068));
  DFRQX1 prev_load_request_reg(.C (rc_gclk), .D (n_349), .Q
       (prev_load_request));
  DFRQX1 prev_read_request_reg(.C (rc_gclk), .D (n_439), .Q (n_6347));
  DFRQX1 prev_write_request_reg(.C (rc_gclk), .D (n_440), .Q (n_6348));
  DFRQX1 \program_counter_reg[0] (.C (rc_gclk_205490), .D (n_432), .Q
       (program_counter[0]));
  DFRQX1 \program_counter_reg[1] (.C (rc_gclk_205490), .D (n_438), .Q
       (program_counter[1]));
  NA2I1X1 g64019(.B (n_1356), .AN (n_971), .Q (n_120));
  NO3I2X1 g52051(.C (n_728), .AN (n_176), .BN (n_6561), .Q (n_119));
  NA2I1X1 g52052(.B (n_872), .AN (n_655), .Q (n_118));
  NA2I1X1 g52054(.B (alu_2nd_operand[20]), .AN (n_4486), .Q (n_116));
  NA2I1X1 g52055(.B (alu_2nd_operand[2]), .AN (n_6628), .Q (n_115));
  NA2I1X1 g52056(.B (n_5542), .AN (n_6373), .Q (n_114));
  AN221X1 g54482(.A (n_270), .B (n_5698), .C (n_135), .D (n_6072), .E
       (n_1546), .Q (n_172));
  AN221X1 g54484(.A (n_270), .B (n_5692), .C (n_135), .D (n_6068), .E
       (n_1529), .Q (n_163));
  AN221X1 g54486(.A (n_270), .B (n_5690), .C (n_135), .D (n_6066), .E
       (n_1532), .Q (n_162));
  AND2X1 g54490(.A (n_119), .B (n_6454), .Q (n_137));
  OA221X1 g54492(.A (n_183), .B (n_273), .C (n_191), .D (n_274), .E
       (n_697), .Q (n_132));
  AN221X1 g54494(.A (n_270), .B (n_5720), .C (n_135), .D (n_6058), .E
       (n_1513), .Q (n_160));
  AN221X1 g54496(.A (n_270), .B (n_5719), .C (n_135), .D (n_6057), .E
       (n_1512), .Q (n_159));
  AN221X1 g54498(.A (n_969), .B (n_1356), .C (n_135), .D (n_6080), .E
       (n_1534), .Q (n_166));
  AND2X2 g54500(.A (n_298), .B (n_6050), .Q (n_130));
  AND2X2 g54502(.A (n_298), .B (n_6051), .Q (n_129));
  INX6 g54504(.A (n_121), .Q (n_123));
  ON21X2 g54506(.A (n_125), .B (n_6048), .C (n_6453), .Q (n_131));
  AND2X1 g54508(.A (n_179), .B (n_4533), .Q (n_127));
  OA221X1 g54510(.A (n_870), .B (n_229), .C (n_869), .D (n_552), .E
       (n_1322), .Q (n_148));
  OA221X1 g54512(.A (n_870), .B (n_222), .C (n_869), .D (n_549), .E
       (n_1319), .Q (n_147));
  OA221X1 g54514(.A (n_870), .B (n_217), .C (n_869), .D (n_557), .E
       (n_1318), .Q (n_146));
  OA221X1 g54516(.A (n_870), .B (n_213), .C (n_869), .D (n_558), .E
       (n_1310), .Q (n_145));
  OA22X1 g54518(.A (n_822), .B (n_964), .C (n_808), .D (n_981), .Q
       (n_140));
  OA221X1 g54520(.A (n_579), .B (n_826), .C (n_572), .D (n_798), .E
       (n_1347), .Q (n_143));
  AND2X2 g54522(.A (n_6453), .B (n_6049), .Q (n_125));
  AND2X2 g54524(.A (n_6048), .B (n_6453), .Q (n_126));
  INX1 g54526(.A (alu_2nd_operand[2]), .Q (n_124));
  AND2X1 g54528(.A (alu_2nd_operand[1]), .B (n_4533), .Q (n_128));
  NO2I1X2 g54530(.B (n_130), .AN (n_568), .Q (n_117));
  INX1 g54532(.A (n_869), .Q (n_133));
  INX1 g54534(.A (n_137), .Q (n_136));
  INX1 g54536(.A (n_870), .Q (n_134));
  OA221X1 g54538(.A (n_869), .B (n_547), .C (n_118), .D (n_790), .E
       (n_1380), .Q (n_150));
  OA221X1 g54540(.A (n_869), .B (n_544), .C (n_118), .D (n_875), .E
       (n_1381), .Q (n_149));
  OA22X1 g54542(.A (n_143), .B (n_871), .C (n_1359), .D (n_977), .Q
       (n_151));
  OA22X1 g54544(.A (n_815), .B (n_973), .C (n_883), .D (n_960), .Q
       (n_138));
  OA22X1 g54546(.A (n_814), .B (n_973), .C (n_879), .D (n_960), .Q
       (n_139));
  OA221X1 g54548(.A (n_960), .B (n_842), .C (n_973), .D (n_805), .E
       (n_1341), .Q (n_142));
  OA221X1 g54550(.A (n_960), .B (n_809), .C (n_958), .D (n_815), .E
       (n_1492), .Q (n_152));
  OA221X1 g54552(.A (n_958), .B (n_816), .C (n_974), .D (n_809), .E
       (n_138), .Q (n_144));
  OA221X1 g54554(.A (n_974), .B (n_806), .C (n_958), .D (n_823), .E
       (n_139), .Q (n_141));
  AND6X1 g54556(.A (n_1062), .B (n_1454), .C (n_566), .D (n_1459), .E
       (n_797), .F (n_1443), .Q (n_155));
  AN221X1 g54558(.A (n_270), .B (n_5696), .C (n_135), .D (n_6070), .E
       (n_1491), .Q (n_153));
  AN221X1 g54560(.A (n_270), .B (n_5694), .C (n_135), .D (n_6069), .E
       (n_1541), .Q (n_170));
  AN221X1 g54562(.A (n_270), .B (n_5688), .C (n_135), .D (n_6063), .E
       (n_1530), .Q (n_164));
  AN221X1 g54564(.A (n_270), .B (n_5686), .C (n_135), .D (n_6062), .E
       (n_1539), .Q (n_169));
  AN221X1 g54566(.A (n_270), .B (n_5684), .C (n_135), .D (n_6061), .E
       (n_1540), .Q (n_168));
  AN221X1 g54568(.A (n_270), .B (n_5722), .C (n_135), .D (n_6060), .E
       (n_1538), .Q (n_167));
  OA221X1 g54570(.A (n_965), .B (n_1006), .C (n_968), .D (n_1366), .E
       (n_152), .Q (n_154));
  AND2X1 g54571(.A (n_5747), .B (n_121), .Q (n_113));
  AND2X1 g54572(.A (n_5737), .B (n_121), .Q (n_112));
  AND2X1 g54573(.A (n_5734), .B (n_121), .Q (n_111));
  AND2X1 g54574(.A (n_5733), .B (n_121), .Q (n_110));
  AND2X1 g54575(.A (n_5731), .B (n_121), .Q (n_109));
  AND2X1 g54576(.A (n_5729), .B (n_121), .Q (n_108));
  AND2X1 g54577(.A (n_5751), .B (n_121), .Q (n_107));
  AND2X1 g54578(.A (n_5750), .B (n_121), .Q (n_106));
  NO2X1 g54581(.A (n_205), .B (n_123), .Q (n_105));
  AND2X1 g54583(.A (n_5748), .B (n_122), .Q (n_104));
  AND2X1 g54585(.A (n_5746), .B (n_122), .Q (n_103));
  AND2X1 g54587(.A (n_4538), .B (n_122), .Q (n_102));
  AND2X1 g54590(.A (n_5743), .B (n_122), .Q (n_101));
  AND2X1 g54593(.A (n_5742), .B (n_122), .Q (n_100));
  AND2X1 g54595(.A (n_5741), .B (n_122), .Q (n_99));
  AND2X1 g54598(.A (n_5740), .B (n_122), .Q (n_98));
  AND2X1 g54600(.A (n_5738), .B (n_122), .Q (n_97));
  AND2X1 g54603(.A (n_5735), .B (n_122), .Q (n_96));
  AND2X1 g54605(.A (n_5732), .B (n_122), .Q (n_95));
  AND2X1 g54607(.A (n_5730), .B (n_122), .Q (n_94));
  AND2X1 g54608(.A (n_6731), .B (n_122), .Q (n_93));
  AND2X1 g54610(.A (n_6730), .B (n_122), .Q (n_92));
  AND2X1 g54611(.A (n_5749), .B (n_122), .Q (n_91));
  AND2X1 g54612(.A (n_4536), .B (n_122), .Q (n_90));
  AND2X1 g54614(.A (n_5739), .B (n_122), .Q (n_89));
  AND2X1 g54616(.A (n_5736), .B (n_122), .Q (n_88));
  AND2X1 g54617(.A (n_5988), .B (n_122), .Q (n_87));
  AND2X1 g54619(.A (n_5987), .B (n_122), .Q (n_86));
  AND2X1 g54620(.A (n_4535), .B (n_122), .Q (n_85));
  AND2X1 g54621(.A (n_5985), .B (n_122), .Q (n_84));
  AND2X1 g54622(.A (n_5729), .B (n_122), .Q (n_83));
  AND2X1 g54623(.A (n_5731), .B (n_122), .Q (n_82));
  AND2X1 g54624(.A (n_5733), .B (n_122), .Q (n_81));
  AND2X1 g54625(.A (n_5734), .B (n_122), .Q (n_80));
  AND2X1 g54626(.A (n_5737), .B (n_122), .Q (n_79));
  NO2X1 g54645(.A (n_1556), .B (n_123), .Q (n_78));
  NO2X1 g54653(.A (n_155), .B (n_123), .Q (n_77));
  NO2X1 g54661(.A (n_153), .B (n_123), .Q (n_76));
  NO2X1 g54673(.A (n_170), .B (n_123), .Q (n_75));
  NO2X1 g54685(.A (n_164), .B (n_123), .Q (n_74));
  NO2X1 g54703(.A (n_169), .B (n_123), .Q (n_73));
  NO2X1 g54725(.A (n_168), .B (n_123), .Q (n_72));
  NO2X1 g54748(.A (n_167), .B (n_123), .Q (n_71));
  NO2X1 g54754(.A (n_165), .B (n_123), .Q (n_70));
  NO2X1 g54780(.A (n_158), .B (n_123), .Q (n_69));
  NO2X1 g54786(.A (n_161), .B (n_123), .Q (n_68));
  NO2X1 g54806(.A (n_1552), .B (n_123), .Q (n_67));
  NO2X1 g54827(.A (n_155), .B (n_123), .Q (n_66));
  NO2X1 g54848(.A (n_153), .B (n_123), .Q (n_65));
  NO2X1 g54871(.A (n_165), .B (n_123), .Q (n_64));
  NO2X2 g54894(.A (n_161), .B (n_123), .Q (n_63));
  NO2X1 g54904(.A (n_1556), .B (n_123), .Q (n_62));
  NO2X1 g54921(.A (n_170), .B (n_123), .Q (n_61));
  NO2X1 g54938(.A (n_164), .B (n_123), .Q (n_60));
  NO2X1 g54949(.A (n_169), .B (n_123), .Q (n_59));
  NO2X1 g54952(.A (n_158), .B (n_123), .Q (n_58));
  NO2X1 g54961(.A (n_1552), .B (n_123), .Q (n_57));
  NO2X1 g54968(.A (n_168), .B (n_123), .Q (n_56));
  NO2X1 g54974(.A (n_167), .B (n_123), .Q (n_55));
  NO2X1 g54986(.A (n_1559), .B (n_123), .Q (n_54));
  NO2X1 g55011(.A (n_172), .B (n_123), .Q (n_53));
  NO2X1 g55023(.A (n_163), .B (n_123), .Q (n_52));
  NO2X1 g55046(.A (n_162), .B (n_123), .Q (n_51));
  NO2X1 g55064(.A (n_171), .B (n_123), .Q (n_50));
  NO2X1 g55080(.A (n_157), .B (n_123), .Q (n_49));
  NO2X1 g55095(.A (n_156), .B (n_123), .Q (n_48));
  NO2X1 g55119(.A (n_1551), .B (n_123), .Q (n_47));
  NO2X1 g55123(.A (n_172), .B (n_123), .Q (n_46));
  NO2X1 g55137(.A (n_156), .B (n_123), .Q (n_45));
  NO2X1 g55154(.A (n_1559), .B (n_123), .Q (n_44));
  NO2X1 g55171(.A (n_163), .B (n_123), .Q (n_43));
  NO2X1 g55184(.A (n_157), .B (n_123), .Q (n_42));
  NO2X1 g55195(.A (n_171), .B (n_123), .Q (n_41));
  NO2X1 g55200(.A (n_1551), .B (n_123), .Q (n_40));
  NO2X1 g55206(.A (n_162), .B (n_123), .Q (n_39));
  NO2X1 g55227(.A (n_1560), .B (n_123), .Q (n_38));
  NO2X1 g55249(.A (n_1549), .B (n_123), .Q (n_37));
  NO2X1 g55267(.A (n_160), .B (n_123), .Q (n_36));
  NO2X1 g55274(.A (n_159), .B (n_123), .Q (n_35));
  NO2X1 g55297(.A (n_1553), .B (n_123), .Q (n_34));
  NO2X1 g55318(.A (n_166), .B (n_123), .Q (n_33));
  NO2X1 g55325(.A (n_1549), .B (n_123), .Q (n_32));
  NO2X1 g55347(.A (n_159), .B (n_123), .Q (n_31));
  NO2X1 g55353(.A (n_1553), .B (n_123), .Q (n_30));
  NO2X1 g55361(.A (n_166), .B (n_123), .Q (n_29));
  NO2X1 g55369(.A (n_1560), .B (n_123), .Q (n_28));
  NO2X1 g55380(.A (n_160), .B (n_123), .Q (n_27));
  NO2X1 g55399(.A (n_1563), .B (n_123), .Q (n_26));
  NO2X1 g55423(.A (n_1555), .B (n_123), .Q (n_25));
  NO2X1 g55432(.A (n_1554), .B (n_123), .Q (n_24));
  NO2X1 g55457(.A (n_1557), .B (n_123), .Q (n_23));
  NO2X1 g55477(.A (n_1554), .B (n_123), .Q (n_22));
  NO2X1 g55487(.A (n_1563), .B (n_123), .Q (n_21));
  NO2X1 g55491(.A (n_1557), .B (n_123), .Q (n_20));
  NO2X1 g55496(.A (n_1555), .B (n_123), .Q (n_19));
  NO2X1 g55503(.A (n_1550), .B (n_123), .Q (n_18));
  NO2X1 g55522(.A (n_1558), .B (n_123), .Q (n_17));
  NO2X1 g55532(.A (n_1558), .B (n_123), .Q (n_16));
  NO2X1 g55554(.A (n_1550), .B (n_123), .Q (n_15));
  AND2X1 g55556(.A (n_119), .B (n_6459), .Q (n_135));
  INX2 g55558(.A (n_123), .Q (n_122));
  AN221X1 g55560(.A (n_270), .B (n_5717), .C (n_135), .D (n_6055), .E
       (n_1547), .Q (n_171));
  AN221X1 g55562(.A (n_270), .B (n_5715), .C (n_135), .D (n_6054), .E
       (n_1515), .Q (n_157));
  AN221X1 g55564(.A (n_270), .B (n_5704), .C (n_135), .D (n_6053), .E
       (n_1508), .Q (n_156));
  AN221X1 g55566(.A (n_270), .B (n_5721), .C (n_135), .D (n_6059), .E
       (n_1531), .Q (n_165));
  AN221X1 g55568(.A (n_270), .B (n_5718), .C (n_135), .D (n_6056), .E
       (n_1514), .Q (n_158));
  AN221X1 g55570(.A (n_270), .B (n_5682), .C (n_135), .D (n_6052), .E
       (n_1511), .Q (n_161));
  OR5X1 g28606(.A (n_13), .B (n_6506), .C (n_6505), .D (n_6503), .E
       (n_6504), .Q (n_14));
  OR6X1 g28608(.A (n_6508), .B (n_6514), .C (n_6510), .D (n_6516), .E
       (n_6512), .F (n_6756), .Q (n_13));
  NO3X1 g28609(.A (n_11), .B (n_6509), .C (n_6512), .Q (n_12));
  OR5X1 g28610(.A (n_6508), .B (n_6513), .C (n_6516), .D (n_6), .E
       (n_6517), .Q (n_11));
  OR6X1 g28613(.A (n_4), .B (n_6514), .C (n_6515), .D (n_6516), .E
       (n_6503), .F (n_2), .Q (n_10));
  OR5X1 g28614(.A (n_4), .B (n_6505), .C (n_7), .D (n_6513), .E
       (n_6510), .Q (n_9));
  OR3X1 g28616(.A (n_6512), .B (n_6511), .C (n_3), .Q (n_7));
  NA6I4X1 g28617(.E (take_trap_39145), .F (n_6238), .AN (n_6519), .BN
       (n_6218), .CN (n_6216), .DN (n_6520), .Q (n_6));
  AN211X1 g28618(.A (n_6217), .B (n_6238), .C (n_3), .D (n_6519), .Q
       (n_5));
  OR4X1 g28619(.A (n_6506), .B (n_6507), .C (n_6508), .D (n_6509), .Q
       (n_4));
  NA2I1X1 g28620(.B (n_1), .AN (n_6517), .Q (n_2));
  NO3I1X1 g28621(.B (n_6596), .C (n_0), .AN (n_5724), .Q (n_3));
  ON21X1 g28622(.A (n_6216), .B (n_6215), .C (n_6238), .Q (n_1));
  NA2X1 g28623(.A (n_6460), .B (n_6238), .Q (n_0));
  EN2X0 add_464_21_g975(.A (add_464_21_n_628), .B (add_464_21_n_803),
       .Q (n_6139));
  EN2X0 add_464_21_g976(.A (add_464_21_n_598), .B (add_464_21_n_802),
       .Q (n_6131));
  EN2X0 add_464_21_g977(.A (add_464_21_n_600), .B (add_464_21_n_816),
       .Q (n_6133));
  EN2X0 add_464_21_g978(.A (add_464_21_n_607), .B (add_464_21_n_813),
       .Q (n_6129));
  EN2X0 add_464_21_g979(.A (add_464_21_n_613), .B (add_464_21_n_809),
       .Q (n_6135));
  EN2X0 add_464_21_g980(.A (add_464_21_n_614), .B (add_464_21_n_810),
       .Q (n_6137));
  EN2X0 add_464_21_g981(.A (add_464_21_n_603), .B (add_464_21_n_815),
       .Q (n_6127));
  EN2X0 add_464_21_g982(.A (add_464_21_n_623), .B (add_464_21_n_789),
       .Q (n_6149));
  EN2X0 add_464_21_g983(.A (add_464_21_n_624), .B (add_464_21_n_808),
       .Q (n_6143));
  EN2X0 add_464_21_g984(.A (add_464_21_n_618), .B (add_464_21_n_773),
       .Q (n_6145));
  EN2X0 add_464_21_g985(.A (add_464_21_n_620), .B (add_464_21_n_782),
       .Q (n_6147));
  EN2X0 add_464_21_g986(.A (add_464_21_n_631), .B (add_464_21_n_805),
       .Q (n_6141));
  EN2X0 add_464_21_g988(.A (add_464_21_n_616), .B (add_464_21_n_792),
       .Q (n_6123));
  EN2X0 add_464_21_g989(.A (add_464_21_n_626), .B (add_464_21_n_763),
       .Q (n_6125));
  EN2X0 add_464_21_g990(.A (add_464_21_n_641), .B (add_464_21_n_783),
       .Q (n_6151));
  AN321X1 add_464_21_g991(.A (add_464_21_n_799), .B (add_464_21_n_712),
       .C (add_464_21_n_640), .D (add_464_21_n_799), .E
       (add_464_21_n_691), .F (add_464_21_n_744), .Q
       (add_464_21_n_598));
  ON321X1 add_464_21_g992(.A (add_464_21_n_916), .B (add_464_21_n_711),
       .C (add_464_21_n_641), .D (add_464_21_n_916), .E
       (add_464_21_n_690), .F (add_464_21_n_910), .Q
       (add_464_21_n_600));
  ON321X1 add_464_21_g993(.A (add_464_21_n_746), .B (add_464_21_n_711),
       .C (add_464_21_n_641), .D (add_464_21_n_746), .E
       (add_464_21_n_690), .F (add_464_21_n_709), .Q
       (add_464_21_n_603));
  AN31X1 add_464_21_g994(.A (add_464_21_n_740), .B (add_464_21_n_712),
       .C (add_464_21_n_640), .D (add_464_21_n_676), .Q
       (add_464_21_n_607));
  AN321X1 add_464_21_g995(.A (add_464_21_n_714), .B (add_464_21_n_712),
       .C (add_464_21_n_640), .D (add_464_21_n_714), .E
       (add_464_21_n_691), .F (add_464_21_n_695), .Q
       (add_464_21_n_610));
  AN21X1 add_464_21_g996(.A (add_464_21_n_640), .B (add_464_21_n_712),
       .C (add_464_21_n_691), .Q (add_464_21_n_613));
  AN31X1 add_464_21_g997(.A (add_464_21_n_742), .B (add_464_21_n_728),
       .C (add_464_21_n_640), .D (add_464_21_n_687), .Q
       (add_464_21_n_614));
  EN2X0 add_464_21_g998(.A (add_464_21_n_639), .B (add_464_21_n_771),
       .Q (n_6153));
  ON321X1 add_464_21_g999(.A (add_464_21_n_716), .B (add_464_21_n_711),
       .C (add_464_21_n_641), .D (add_464_21_n_716), .E
       (add_464_21_n_690), .F (add_464_21_n_697), .Q
       (add_464_21_n_616));
  AN321X1 add_464_21_g1000(.A (add_464_21_n_860), .B
       (add_464_21_n_759), .C (add_464_21_n_640), .D
       (add_464_21_n_860), .E (add_464_21_n_727), .F
       (add_464_21_n_852), .Q (add_464_21_n_618));
  AN21X1 add_464_21_g1001(.A (add_464_21_n_640), .B (add_464_21_n_759),
       .C (add_464_21_n_727), .Q (add_464_21_n_620));
  ON21X1 add_464_21_g1002(.A (add_464_21_n_641), .B (add_464_21_n_845),
       .C (add_464_21_n_850), .Q (add_464_21_n_623));
  AN21X1 add_464_21_g1003(.A (add_464_21_n_640), .B (add_464_21_n_728),
       .C (add_464_21_n_702), .Q (add_464_21_n_624));
  AN321X1 add_464_21_g1004(.A (add_464_21_n_718), .B
       (add_464_21_n_712), .C (add_464_21_n_640), .D
       (add_464_21_n_718), .E (add_464_21_n_691), .F
       (add_464_21_n_699), .Q (add_464_21_n_626));
  AN321X1 add_464_21_g1005(.A (add_464_21_n_800), .B
       (add_464_21_n_728), .C (add_464_21_n_640), .D
       (add_464_21_n_800), .E (add_464_21_n_702), .F
       (add_464_21_n_743), .Q (add_464_21_n_628));
  ON321X1 add_464_21_g1006(.A (add_464_21_n_920), .B
       (add_464_21_n_729), .C (add_464_21_n_641), .D
       (add_464_21_n_920), .E (add_464_21_n_703), .F
       (add_464_21_n_897), .Q (add_464_21_n_631));
  EN2X0 add_464_21_g1007(.A (add_464_21_n_644), .B (add_464_21_n_780),
       .Q (n_6159));
  EN2X0 add_464_21_g1008(.A (add_464_21_n_662), .B (add_464_21_n_824),
       .Q (n_6165));
  EN2X0 add_464_21_g1009(.A (add_464_21_n_652), .B (add_464_21_n_786),
       .Q (n_6157));
  EN2X0 add_464_21_g1010(.A (add_464_21_n_650), .B (add_464_21_n_785),
       .Q (n_6155));
  EN2X0 add_464_21_g1011(.A (add_464_21_n_656), .B (add_464_21_n_777),
       .Q (n_6161));
  EN2X0 add_464_21_g1012(.A (add_464_21_n_659), .B (add_464_21_n_829),
       .Q (n_6163));
  AN21X1 add_464_21_g1013(.A (add_464_21_n_663), .B (add_464_21_n_722),
       .C (add_464_21_n_692), .Q (add_464_21_n_639));
  INX1 add_464_21_g1014(.A (add_464_21_n_640), .Q (add_464_21_n_641));
  AO221X1 add_464_21_g1015(.A (add_464_21_n_721), .B
       (add_464_21_n_663), .C (add_464_21_n_707), .D
       (add_464_21_n_721), .E (add_464_21_n_705), .Q
       (add_464_21_n_640));
  NO2X1 add_464_21_g1016(.A (add_464_21_n_663), .B (add_464_21_n_707),
       .Q (add_464_21_n_644));
  EN2X1 add_464_21_g1017(.A (add_464_21_n_673), .B (add_464_21_n_819),
       .Q (n_6171));
  EN2X0 add_464_21_g1018(.A (add_464_21_n_674), .B (add_464_21_n_827),
       .Q (n_6173));
  EN2X1 add_464_21_g1019(.A (add_464_21_n_665), .B (add_464_21_n_830),
       .Q (n_6167));
  EN2X1 add_464_21_g1020(.A (add_464_21_n_669), .B (add_464_21_n_821),
       .Q (n_6169));
  AN321X1 add_464_21_g1021(.A (add_464_21_n_762), .B
       (add_464_21_n_726), .C (add_464_21_n_666), .D
       (add_464_21_n_762), .E (add_464_21_n_707), .F
       (add_464_21_n_724), .Q (add_464_21_n_650));
  AO321X1 add_464_21_g1022(.A (add_464_21_n_859), .B
       (add_464_21_n_726), .C (add_464_21_n_666), .D
       (add_464_21_n_859), .E (add_464_21_n_707), .F
       (add_464_21_n_855), .Q (add_464_21_n_652));
  ON321X1 add_464_21_g1023(.A (add_464_21_n_915), .B
       (add_464_21_n_798), .C (add_464_21_n_665), .D
       (add_464_21_n_915), .E (add_464_21_n_745), .F
       (add_464_21_n_907), .Q (add_464_21_n_656));
  OA21X1 add_464_21_g1024(.A (add_464_21_n_665), .B (add_464_21_n_798),
       .C (add_464_21_n_745), .Q (add_464_21_n_659));
  ON21X1 add_464_21_g1025(.A (add_464_21_n_665), .B (add_464_21_n_902),
       .C (add_464_21_n_914), .Q (add_464_21_n_662));
  AND2X1 add_464_21_g1026(.A (add_464_21_n_666), .B (add_464_21_n_726),
       .Q (add_464_21_n_663));
  EN2X1 add_464_21_g1027(.A (add_464_21_n_680), .B (add_464_21_n_768),
       .Q (n_6175));
  INX1 add_464_21_g1028(.A (add_464_21_n_665), .Q (add_464_21_n_666));
  AN321X1 add_464_21_g1029(.A (add_464_21_n_797), .B
       (add_464_21_n_761), .C (add_464_21_n_680), .D
       (add_464_21_n_797), .E (add_464_21_n_725), .F
       (add_464_21_n_748), .Q (add_464_21_n_665));
  AN321X1 add_464_21_g1030(.A (add_464_21_n_917), .B
       (add_464_21_n_761), .C (add_464_21_n_680), .D
       (add_464_21_n_917), .E (add_464_21_n_725), .F
       (add_464_21_n_909), .Q (add_464_21_n_669));
  AN21X1 add_464_21_g1031(.A (add_464_21_n_680), .B (add_464_21_n_761),
       .C (add_464_21_n_725), .Q (add_464_21_n_673));
  ON21X1 add_464_21_g1032(.A (add_464_21_n_681), .B (add_464_21_n_847),
       .C (add_464_21_n_857), .Q (add_464_21_n_674));
  EN2X1 add_464_21_g1033(.A (add_464_21_n_684), .B (add_464_21_n_775),
       .Q (n_6177));
  AO221X1 add_464_21_g1034(.A (add_464_21_n_740), .B
       (add_464_21_n_691), .C (add_464_21_n_919), .D
       (add_464_21_n_744), .E (add_464_21_n_898), .Q
       (add_464_21_n_676));
  EN2X1 add_464_21_g1035(.A (add_464_21_n_700), .B (add_464_21_n_770),
       .Q (n_6179));
  INX1 add_464_21_g1036(.A (add_464_21_n_680), .Q (add_464_21_n_681));
  AO321X1 add_464_21_g1037(.A (add_464_21_n_848), .B
       (add_464_21_n_849), .C (add_464_21_n_700), .D
       (add_464_21_n_843), .E (add_464_21_n_849), .F
       (add_464_21_n_832), .Q (add_464_21_n_680));
  AN21X1 add_464_21_g1038(.A (add_464_21_n_700), .B (add_464_21_n_848),
       .C (add_464_21_n_843), .Q (add_464_21_n_684));
  AO221X1 add_464_21_g1039(.A (add_464_21_n_742), .B
       (add_464_21_n_702), .C (add_464_21_n_918), .D
       (add_464_21_n_743), .E (add_464_21_n_912), .Q
       (add_464_21_n_687));
  INX1 add_464_21_g1040(.A (add_464_21_n_690), .Q (add_464_21_n_691));
  AN221X1 add_464_21_g1041(.A (add_464_21_n_796), .B
       (add_464_21_n_743), .C (add_464_21_n_720), .D
       (add_464_21_n_702), .E (add_464_21_n_747), .Q
       (add_464_21_n_690));
  AO221X1 add_464_21_g1042(.A (add_464_21_n_722), .B
       (add_464_21_n_707), .C (add_464_21_n_858), .D
       (add_464_21_n_724), .E (add_464_21_n_840), .Q
       (add_464_21_n_692));
  ON221X1 add_464_21_g1043(.A (add_464_21_n_723), .B
       (add_464_21_n_709), .C (add_464_21_n_853), .D
       (add_464_21_n_741), .E (add_464_21_n_835), .Q
       (add_464_21_n_695));
  OA21X1 add_464_21_g1044(.A (add_464_21_n_709), .B (add_464_21_n_760),
       .C (add_464_21_n_741), .Q (add_464_21_n_697));
  ON21X1 add_464_21_g1045(.A (add_464_21_n_709), .B (add_464_21_n_861),
       .C (add_464_21_n_856), .Q (add_464_21_n_699));
  FAX1 add_464_21_g1046(.A (program_counter[1]), .B (n_6716), .CI
       (add_464_21_n_731), .S (n_6181), .CO (add_464_21_n_700));
  INX1 add_464_21_g1047(.A (add_464_21_n_703), .Q (add_464_21_n_702));
  AN221X1 add_464_21_g1048(.A (add_464_21_n_852), .B
       (add_464_21_n_844), .C (add_464_21_n_756), .D
       (add_464_21_n_727), .E (add_464_21_n_836), .Q
       (add_464_21_n_703));
  AO221X1 add_464_21_g1049(.A (add_464_21_n_757), .B
       (add_464_21_n_724), .C (add_464_21_n_840), .D
       (add_464_21_n_846), .E (add_464_21_n_839), .Q
       (add_464_21_n_705));
  ON221X1 add_464_21_g1050(.A (add_464_21_n_745), .B
       (add_464_21_n_758), .C (add_464_21_n_907), .D
       (add_464_21_n_851), .E (add_464_21_n_837), .Q
       (add_464_21_n_707));
  AN221X1 add_464_21_g1051(.A (add_464_21_n_898), .B
       (add_464_21_n_906), .C (add_464_21_n_795), .D
       (add_464_21_n_744), .E (add_464_21_n_891), .Q
       (add_464_21_n_709));
  INX1 add_464_21_g1052(.A (add_464_21_n_711), .Q (add_464_21_n_712));
  NA2X1 add_464_21_g1053(.A (add_464_21_n_728), .B (add_464_21_n_720),
       .Q (add_464_21_n_711));
  NO2X1 add_464_21_g1054(.A (add_464_21_n_746), .B (add_464_21_n_723),
       .Q (add_464_21_n_714));
  OR2X1 add_464_21_g1055(.A (add_464_21_n_746), .B (add_464_21_n_760),
       .Q (add_464_21_n_716));
  NO2X1 add_464_21_g1056(.A (add_464_21_n_746), .B (add_464_21_n_861),
       .Q (add_464_21_n_718));
  INX1 add_464_21_g1057(.A (add_464_21_n_728), .Q (add_464_21_n_729));
  HAX1 add_464_21_g1058(.A (n_6014), .B (program_counter[0]), .S
       (n_6183), .CO (add_464_21_n_731));
  AND2X1 add_464_21_g1059(.A (add_464_21_n_796), .B (add_464_21_n_800),
       .Q (add_464_21_n_720));
  AND2X1 add_464_21_g1060(.A (add_464_21_n_757), .B (add_464_21_n_762),
       .Q (add_464_21_n_721));
  AND2X1 add_464_21_g1061(.A (add_464_21_n_762), .B (add_464_21_n_858),
       .Q (add_464_21_n_722));
  OR2X1 add_464_21_g1062(.A (add_464_21_n_760), .B (add_464_21_n_853),
       .Q (add_464_21_n_723));
  ON21X1 add_464_21_g1063(.A (add_464_21_n_854), .B (add_464_21_n_841),
       .C (add_464_21_n_834), .Q (add_464_21_n_724));
  ON21X1 add_464_21_g1064(.A (add_464_21_n_857), .B (add_464_21_n_901),
       .C (add_464_21_n_895), .Q (add_464_21_n_725));
  NO2X1 add_464_21_g1065(.A (add_464_21_n_758), .B (add_464_21_n_798),
       .Q (add_464_21_n_726));
  ON21X1 add_464_21_g1066(.A (add_464_21_n_850), .B (add_464_21_n_842),
       .C (add_464_21_n_838), .Q (add_464_21_n_727));
  AND2X1 add_464_21_g1067(.A (add_464_21_n_756), .B (add_464_21_n_759),
       .Q (add_464_21_n_728));
  ON21X1 add_464_21_g1068(.A (add_464_21_n_911), .B (add_464_21_n_899),
       .C (add_464_21_n_893), .Q (add_464_21_n_747));
  ON21X1 add_464_21_g1069(.A (add_464_21_n_900), .B (add_464_21_n_908),
       .C (add_464_21_n_894), .Q (add_464_21_n_748));
  AND2X1 add_464_21_g1070(.A (add_464_21_n_799), .B (add_464_21_n_919),
       .Q (add_464_21_n_740));
  OA21X1 add_464_21_g1071(.A (add_464_21_n_856), .B (add_464_21_n_904),
       .C (add_464_21_n_833), .Q (add_464_21_n_741));
  AND2X1 add_464_21_g1072(.A (add_464_21_n_800), .B (add_464_21_n_918),
       .Q (add_464_21_n_742));
  ON21X1 add_464_21_g1073(.A (add_464_21_n_897), .B (add_464_21_n_903),
       .C (add_464_21_n_896), .Q (add_464_21_n_743));
  ON21X1 add_464_21_g1074(.A (add_464_21_n_910), .B (add_464_21_n_913),
       .C (add_464_21_n_892), .Q (add_464_21_n_744));
  OA21X1 add_464_21_g1075(.A (add_464_21_n_914), .B (add_464_21_n_905),
       .C (add_464_21_n_890), .Q (add_464_21_n_745));
  NA2X1 add_464_21_g1076(.A (add_464_21_n_795), .B (add_464_21_n_799),
       .Q (add_464_21_n_746));
  NO2I1X1 add_464_21_g1077(.B (add_464_21_n_904), .AN
       (add_464_21_n_833), .Q (add_464_21_n_763));
  AND2X1 add_464_21_g1078(.A (add_464_21_n_844), .B (add_464_21_n_860),
       .Q (add_464_21_n_756));
  AND2X1 add_464_21_g1079(.A (add_464_21_n_846), .B (add_464_21_n_858),
       .Q (add_464_21_n_757));
  NA2I1X1 add_464_21_g1080(.B (add_464_21_n_857), .AN
       (add_464_21_n_847), .Q (add_464_21_n_768));
  NA2I1X1 add_464_21_g1081(.B (add_464_21_n_848), .AN
       (add_464_21_n_843), .Q (add_464_21_n_770));
  NO2I1X1 add_464_21_g1082(.B (add_464_21_n_839), .AN
       (add_464_21_n_846), .Q (add_464_21_n_771));
  NO2I1X1 add_464_21_g1083(.B (add_464_21_n_836), .AN
       (add_464_21_n_844), .Q (add_464_21_n_773));
  NO2I1X1 add_464_21_g1084(.B (add_464_21_n_832), .AN
       (add_464_21_n_849), .Q (add_464_21_n_775));
  NA2I1X1 add_464_21_g1085(.B (add_464_21_n_837), .AN
       (add_464_21_n_851), .Q (add_464_21_n_777));
  AND2X1 add_464_21_g1086(.A (add_464_21_n_859), .B (add_464_21_n_854),
       .Q (add_464_21_n_780));
  NO2I1X1 add_464_21_g1087(.B (add_464_21_n_852), .AN
       (add_464_21_n_860), .Q (add_464_21_n_782));
  NO2I1X1 add_464_21_g1088(.B (add_464_21_n_845), .AN
       (add_464_21_n_850), .Q (add_464_21_n_783));
  NO2I1X1 add_464_21_g1089(.B (add_464_21_n_840), .AN
       (add_464_21_n_858), .Q (add_464_21_n_785));
  NA2I1X1 add_464_21_g1090(.B (add_464_21_n_834), .AN
       (add_464_21_n_841), .Q (add_464_21_n_786));
  NA2I1X1 add_464_21_g1091(.B (add_464_21_n_838), .AN
       (add_464_21_n_842), .Q (add_464_21_n_789));
  NA2I1X1 add_464_21_g1092(.B (add_464_21_n_835), .AN
       (add_464_21_n_853), .Q (add_464_21_n_792));
  OR2X1 add_464_21_g1093(.A (add_464_21_n_851), .B (add_464_21_n_915),
       .Q (add_464_21_n_758));
  NO2X1 add_464_21_g1094(.A (add_464_21_n_845), .B (add_464_21_n_842),
       .Q (add_464_21_n_759));
  OR2X1 add_464_21_g1095(.A (add_464_21_n_904), .B (add_464_21_n_861),
       .Q (add_464_21_n_760));
  NO2X1 add_464_21_g1096(.A (add_464_21_n_847), .B (add_464_21_n_901),
       .Q (add_464_21_n_761));
  NO2I1X1 add_464_21_g1097(.B (add_464_21_n_841), .AN
       (add_464_21_n_859), .Q (add_464_21_n_762));
  AND2X1 add_464_21_g1098(.A (add_464_21_n_906), .B (add_464_21_n_919),
       .Q (add_464_21_n_795));
  NO2I1X1 add_464_21_g1099(.B (add_464_21_n_898), .AN
       (add_464_21_n_919), .Q (add_464_21_n_802));
  AND2X1 add_464_21_g1100(.A (add_464_21_n_918), .B (add_464_21_n_911),
       .Q (add_464_21_n_803));
  NA2I1X1 add_464_21_g1101(.B (add_464_21_n_896), .AN
       (add_464_21_n_903), .Q (add_464_21_n_805));
  NO2I1X1 add_464_21_g1102(.B (add_464_21_n_920), .AN
       (add_464_21_n_897), .Q (add_464_21_n_808));
  NO2I1X1 add_464_21_g1103(.B (add_464_21_n_916), .AN
       (add_464_21_n_910), .Q (add_464_21_n_809));
  NO2I1X1 add_464_21_g1104(.B (add_464_21_n_899), .AN
       (add_464_21_n_893), .Q (add_464_21_n_810));
  NO2I1X1 add_464_21_g1105(.B (add_464_21_n_891), .AN
       (add_464_21_n_906), .Q (add_464_21_n_813));
  NA2I1X1 add_464_21_g1106(.B (add_464_21_n_856), .AN
       (add_464_21_n_861), .Q (add_464_21_n_815));
  NA2I1X1 add_464_21_g1107(.B (add_464_21_n_892), .AN
       (add_464_21_n_913), .Q (add_464_21_n_816));
  AND2X1 add_464_21_g1108(.A (add_464_21_n_917), .B (add_464_21_n_908),
       .Q (add_464_21_n_819));
  NO2I1X1 add_464_21_g1109(.B (add_464_21_n_899), .AN
       (add_464_21_n_918), .Q (add_464_21_n_796));
  NO2I1X1 add_464_21_g1110(.B (add_464_21_n_900), .AN
       (add_464_21_n_894), .Q (add_464_21_n_821));
  NO2I1X1 add_464_21_g1111(.B (add_464_21_n_900), .AN
       (add_464_21_n_917), .Q (add_464_21_n_797));
  NA2I1X1 add_464_21_g1112(.B (add_464_21_n_890), .AN
       (add_464_21_n_905), .Q (add_464_21_n_824));
  NA2I1X1 add_464_21_g1113(.B (add_464_21_n_895), .AN
       (add_464_21_n_901), .Q (add_464_21_n_827));
  NO2I1X1 add_464_21_g1114(.B (add_464_21_n_915), .AN
       (add_464_21_n_907), .Q (add_464_21_n_829));
  NO2I1X1 add_464_21_g1115(.B (add_464_21_n_902), .AN
       (add_464_21_n_914), .Q (add_464_21_n_830));
  OR2X1 add_464_21_g1116(.A (add_464_21_n_902), .B (add_464_21_n_905),
       .Q (add_464_21_n_798));
  NO2X1 add_464_21_g1117(.A (add_464_21_n_916), .B (add_464_21_n_913),
       .Q (add_464_21_n_799));
  NO2X1 add_464_21_g1118(.A (add_464_21_n_920), .B (add_464_21_n_903),
       .Q (add_464_21_n_800));
  INX1 add_464_21_g1119(.A (add_464_21_n_854), .Q (add_464_21_n_855));
  AND2X1 add_464_21_g1120(.A (n_6010), .B (program_counter[3]), .Q
       (add_464_21_n_832));
  NA2X1 add_464_21_g1121(.A (n_5994), .B (program_counter[29]), .Q
       (add_464_21_n_833));
  NA2X1 add_464_21_g1122(.A (n_6007), .B (program_counter[13]), .Q
       (add_464_21_n_834));
  NA2X1 add_464_21_g1123(.A (n_5993), .B (program_counter[30]), .Q
       (add_464_21_n_835));
  AND2X1 add_464_21_g1124(.A (n_6001), .B (program_counter[19]), .Q
       (add_464_21_n_836));
  NA2X1 add_464_21_g1125(.A (n_6013), .B (program_counter[11]), .Q
       (add_464_21_n_837));
  NA2X1 add_464_21_g1126(.A (n_6003), .B (program_counter[17]), .Q
       (add_464_21_n_838));
  AND2X1 add_464_21_g1127(.A (n_6005), .B (program_counter[15]), .Q
       (add_464_21_n_839));
  AND2X1 add_464_21_g1128(.A (n_6006), .B (program_counter[14]), .Q
       (add_464_21_n_840));
  NO2X1 add_464_21_g1129(.A (n_6007), .B (program_counter[13]), .Q
       (add_464_21_n_841));
  NO2X1 add_464_21_g1130(.A (n_6003), .B (program_counter[17]), .Q
       (add_464_21_n_842));
  AND2X1 add_464_21_g1131(.A (n_6011), .B (program_counter[2]), .Q
       (add_464_21_n_843));
  OR2X1 add_464_21_g1132(.A (n_6001), .B (program_counter[19]), .Q
       (add_464_21_n_844));
  NO2X1 add_464_21_g1133(.A (n_6004), .B (program_counter[16]), .Q
       (add_464_21_n_845));
  OR2X1 add_464_21_g1134(.A (n_6005), .B (program_counter[15]), .Q
       (add_464_21_n_846));
  NO2X1 add_464_21_g1135(.A (n_6717), .B (program_counter[4]), .Q
       (add_464_21_n_847));
  OR2X1 add_464_21_g1136(.A (n_6011), .B (program_counter[2]), .Q
       (add_464_21_n_848));
  OR2X1 add_464_21_g1137(.A (n_6010), .B (program_counter[3]), .Q
       (add_464_21_n_849));
  NA2X1 add_464_21_g1138(.A (n_6004), .B (program_counter[16]), .Q
       (add_464_21_n_850));
  NO2X1 add_464_21_g1139(.A (n_6013), .B (program_counter[11]), .Q
       (add_464_21_n_851));
  AND2X1 add_464_21_g1140(.A (n_6002), .B (program_counter[18]), .Q
       (add_464_21_n_852));
  NO2X1 add_464_21_g1141(.A (n_5993), .B (program_counter[30]), .Q
       (add_464_21_n_853));
  NA2X1 add_464_21_g1142(.A (n_6008), .B (program_counter[12]), .Q
       (add_464_21_n_854));
  NA2X1 add_464_21_g1143(.A (n_5995), .B (program_counter[28]), .Q
       (add_464_21_n_856));
  NA2X1 add_464_21_g1144(.A (n_6717), .B (program_counter[4]), .Q
       (add_464_21_n_857));
  OR2X1 add_464_21_g1145(.A (n_6006), .B (program_counter[14]), .Q
       (add_464_21_n_858));
  OR2X1 add_464_21_g1146(.A (n_6008), .B (program_counter[12]), .Q
       (add_464_21_n_859));
  OR2X1 add_464_21_g1147(.A (n_6002), .B (program_counter[18]), .Q
       (add_464_21_n_860));
  NO2X1 add_464_21_g1148(.A (n_5995), .B (program_counter[28]), .Q
       (add_464_21_n_861));
  INX1 add_464_21_g1149(.A (add_464_21_n_908), .Q (add_464_21_n_909));
  INX1 add_464_21_g1150(.A (add_464_21_n_911), .Q (add_464_21_n_912));
  NA2X1 add_464_21_g1151(.A (n_6558), .B (program_counter[9]), .Q
       (add_464_21_n_890));
  AND2X1 add_464_21_g1152(.A (n_5996), .B (program_counter[27]), .Q
       (add_464_21_n_891));
  NA2X1 add_464_21_g1153(.A (n_5998), .B (program_counter[25]), .Q
       (add_464_21_n_892));
  NA2X1 add_464_21_g1154(.A (n_6000), .B (program_counter[23]), .Q
       (add_464_21_n_893));
  NA2X1 add_464_21_g1155(.A (n_6556), .B (program_counter[7]), .Q
       (add_464_21_n_894));
  NA2X1 add_464_21_g1156(.A (n_6554), .B (program_counter[5]), .Q
       (add_464_21_n_895));
  NA2X1 add_464_21_g1157(.A (n_6015), .B (program_counter[21]), .Q
       (add_464_21_n_896));
  NA2X1 add_464_21_g1158(.A (n_5992), .B (program_counter[20]), .Q
       (add_464_21_n_897));
  AND2X1 add_464_21_g1159(.A (n_5997), .B (program_counter[26]), .Q
       (add_464_21_n_898));
  NO2X1 add_464_21_g1160(.A (n_6000), .B (program_counter[23]), .Q
       (add_464_21_n_899));
  NO2X1 add_464_21_g1161(.A (n_6556), .B (program_counter[7]), .Q
       (add_464_21_n_900));
  NO2X1 add_464_21_g1162(.A (n_6554), .B (program_counter[5]), .Q
       (add_464_21_n_901));
  NO2X1 add_464_21_g1163(.A (n_6557), .B (program_counter[8]), .Q
       (add_464_21_n_902));
  NO2X1 add_464_21_g1164(.A (n_6015), .B (program_counter[21]), .Q
       (add_464_21_n_903));
  NO2X1 add_464_21_g1165(.A (n_5994), .B (program_counter[29]), .Q
       (add_464_21_n_904));
  NO2X1 add_464_21_g1166(.A (n_6558), .B (program_counter[9]), .Q
       (add_464_21_n_905));
  OR2X1 add_464_21_g1167(.A (n_5996), .B (program_counter[27]), .Q
       (add_464_21_n_906));
  NA2X1 add_464_21_g1168(.A (n_6559), .B (program_counter[10]), .Q
       (add_464_21_n_907));
  NA2X1 add_464_21_g1169(.A (n_6555), .B (program_counter[6]), .Q
       (add_464_21_n_908));
  NA2X1 add_464_21_g1170(.A (n_5999), .B (program_counter[24]), .Q
       (add_464_21_n_910));
  NA2X1 add_464_21_g1171(.A (n_5991), .B (program_counter[22]), .Q
       (add_464_21_n_911));
  NO2X1 add_464_21_g1172(.A (n_5998), .B (program_counter[25]), .Q
       (add_464_21_n_913));
  NA2X1 add_464_21_g1173(.A (n_6557), .B (program_counter[8]), .Q
       (add_464_21_n_914));
  NO2X1 add_464_21_g1174(.A (n_6559), .B (program_counter[10]), .Q
       (add_464_21_n_915));
  NO2X1 add_464_21_g1175(.A (n_5999), .B (program_counter[24]), .Q
       (add_464_21_n_916));
  OR2X1 add_464_21_g1176(.A (n_6555), .B (program_counter[6]), .Q
       (add_464_21_n_917));
  OR2X1 add_464_21_g1177(.A (n_5991), .B (program_counter[22]), .Q
       (add_464_21_n_918));
  OR2X1 add_464_21_g1178(.A (n_5997), .B (program_counter[26]), .Q
       (add_464_21_n_919));
  NO2X1 add_464_21_g1179(.A (n_5992), .B (program_counter[20]), .Q
       (add_464_21_n_920));
  EN3X1 add_464_21_g1181(.A (add_464_21_n_610), .B (n_6560), .C
       (program_counter[31]), .Q (n_6121));
  EN2X0 add_463_14_g969(.A (add_463_14_n_636), .B (add_463_14_n_807),
       .Q (n_6148));
  EN2X0 add_463_14_g970(.A (add_463_14_n_598), .B (add_463_14_n_788),
       .Q (n_6132));
  EN2X0 add_463_14_g971(.A (add_463_14_n_601), .B (add_463_14_n_805),
       .Q (n_6134));
  EN2X0 add_463_14_g972(.A (add_463_14_n_608), .B (add_463_14_n_776),
       .Q (n_6130));
  EN2X0 add_463_14_g973(.A (add_463_14_n_613), .B (add_463_14_n_809),
       .Q (n_6136));
  EN2X0 add_463_14_g974(.A (add_463_14_n_620), .B (add_463_14_n_802),
       .Q (n_6144));
  EN2X0 add_463_14_g975(.A (add_463_14_n_603), .B (add_463_14_n_784),
       .Q (n_6128));
  EN2X0 add_463_14_g976(.A (add_463_14_n_614), .B (add_463_14_n_771),
       .Q (n_6138));
  EN2X0 add_463_14_g977(.A (add_463_14_n_615), .B (add_463_14_n_789),
       .Q (n_6140));
  EN2X0 add_463_14_g978(.A (add_463_14_n_618), .B (add_463_14_n_800),
       .Q (n_6142));
  EN2X0 add_463_14_g979(.A (add_463_14_n_633), .B (add_463_14_n_817),
       .Q (n_6146));
  EN2X0 add_463_14_g980(.A (add_463_14_n_635), .B (add_463_14_n_821),
       .Q (n_6150));
  EN2X0 add_463_14_g982(.A (add_463_14_n_629), .B (add_463_14_n_780),
       .Q (n_6124));
  EN2X0 add_463_14_g983(.A (add_463_14_n_631), .B (add_463_14_n_785),
       .Q (n_6126));
  EN2X0 add_463_14_g984(.A (add_463_14_n_654), .B (add_463_14_n_812),
       .Q (n_6152));
  AN321X1 add_463_14_g985(.A (add_463_14_n_764), .B (add_463_14_n_717),
       .C (add_463_14_n_654), .D (add_463_14_n_764), .E
       (add_463_14_n_695), .F (add_463_14_n_739), .Q
       (add_463_14_n_598));
  ON321X1 add_463_14_g986(.A (add_463_14_n_854), .B (add_463_14_n_716),
       .C (add_463_14_n_655), .D (add_463_14_n_854), .E
       (add_463_14_n_694), .F (add_463_14_n_903), .Q
       (add_463_14_n_601));
  ON321X1 add_463_14_g987(.A (add_463_14_n_727), .B (add_463_14_n_716),
       .C (add_463_14_n_655), .D (add_463_14_n_727), .E
       (add_463_14_n_694), .F (add_463_14_n_698), .Q
       (add_463_14_n_603));
  AN31X1 add_463_14_g988(.A (add_463_14_n_724), .B (add_463_14_n_717),
       .C (add_463_14_n_654), .D (add_463_14_n_673), .Q
       (add_463_14_n_608));
  AN321X1 add_463_14_g989(.A (add_463_14_n_717), .B (add_463_14_n_710),
       .C (add_463_14_n_654), .D (add_463_14_n_710), .E
       (add_463_14_n_695), .F (add_463_14_n_683), .Q
       (add_463_14_n_610));
  AN21X1 add_463_14_g990(.A (add_463_14_n_654), .B (add_463_14_n_717),
       .C (add_463_14_n_695), .Q (add_463_14_n_613));
  AN31X1 add_463_14_g991(.A (add_463_14_n_723), .B (add_463_14_n_725),
       .C (add_463_14_n_654), .D (add_463_14_n_688), .Q
       (add_463_14_n_614));
  AN321X1 add_463_14_g992(.A (add_463_14_n_763), .B (add_463_14_n_725),
       .C (add_463_14_n_654), .D (add_463_14_n_763), .E
       (add_463_14_n_705), .F (add_463_14_n_744), .Q
       (add_463_14_n_615));
  ON321X1 add_463_14_g993(.A (add_463_14_n_851), .B (add_463_14_n_726),
       .C (add_463_14_n_655), .D (add_463_14_n_851), .E
       (add_463_14_n_706), .F (add_463_14_n_887), .Q
       (add_463_14_n_618));
  AN21X1 add_463_14_g994(.A (add_463_14_n_654), .B (add_463_14_n_725),
       .C (add_463_14_n_705), .Q (add_463_14_n_620));
  EN2X0 add_463_14_g995(.A (add_463_14_n_644), .B (add_463_14_n_803),
       .Q (n_6158));
  EN2X0 add_463_14_g996(.A (add_463_14_n_639), .B (add_463_14_n_774),
       .Q (n_6154));
  EN2X0 add_463_14_g997(.A (add_463_14_n_648), .B (add_463_14_n_766),
       .Q (n_6162));
  EN2X0 add_463_14_g998(.A (add_463_14_n_647), .B (add_463_14_n_798),
       .Q (n_6160));
  EN2X0 add_463_14_g999(.A (add_463_14_n_650), .B (add_463_14_n_816),
       .Q (n_6164));
  EN2X0 add_463_14_g1000(.A (add_463_14_n_640), .B (add_463_14_n_791),
       .Q (n_6156));
  EN2X1 add_463_14_g1001(.A (add_463_14_n_653), .B (add_463_14_n_826),
       .Q (n_6166));
  ON321X1 add_463_14_g1002(.A (add_463_14_n_716), .B
       (add_463_14_n_712), .C (add_463_14_n_655), .D
       (add_463_14_n_712), .E (add_463_14_n_694), .F
       (add_463_14_n_685), .Q (add_463_14_n_629));
  AN321X1 add_463_14_g1003(.A (add_463_14_n_714), .B
       (add_463_14_n_717), .C (add_463_14_n_654), .D
       (add_463_14_n_714), .E (add_463_14_n_695), .F
       (add_463_14_n_687), .Q (add_463_14_n_631));
  AN321X1 add_463_14_g1004(.A (add_463_14_n_855), .B
       (add_463_14_n_796), .C (add_463_14_n_654), .D
       (add_463_14_n_855), .E (add_463_14_n_742), .F
       (add_463_14_n_901), .Q (add_463_14_n_633));
  ON21X1 add_463_14_g1005(.A (add_463_14_n_655), .B (add_463_14_n_892),
       .C (add_463_14_n_894), .Q (add_463_14_n_635));
  AN21X1 add_463_14_g1006(.A (add_463_14_n_654), .B (add_463_14_n_796),
       .C (add_463_14_n_742), .Q (add_463_14_n_636));
  AN31X1 add_463_14_g1007(.A (add_463_14_n_719), .B (add_463_14_n_728),
       .C (add_463_14_n_663), .D (add_463_14_n_691), .Q
       (add_463_14_n_639));
  AN321X1 add_463_14_g1008(.A (add_463_14_n_765), .B
       (add_463_14_n_728), .C (add_463_14_n_663), .D
       (add_463_14_n_765), .E (add_463_14_n_708), .F
       (add_463_14_n_740), .Q (add_463_14_n_640));
  AO321X1 add_463_14_g1009(.A (add_463_14_n_852), .B
       (add_463_14_n_728), .C (add_463_14_n_663), .D
       (add_463_14_n_852), .E (add_463_14_n_708), .F
       (add_463_14_n_906), .Q (add_463_14_n_644));
  AO21X1 add_463_14_g1010(.A (add_463_14_n_663), .B (add_463_14_n_728),
       .C (add_463_14_n_708), .Q (add_463_14_n_647));
  AO321X1 add_463_14_g1011(.A (add_463_14_n_853), .B
       (add_463_14_n_795), .C (add_463_14_n_663), .D
       (add_463_14_n_853), .E (add_463_14_n_743), .F
       (add_463_14_n_904), .Q (add_463_14_n_648));
  AN21X1 add_463_14_g1012(.A (add_463_14_n_663), .B (add_463_14_n_795),
       .C (add_463_14_n_743), .Q (add_463_14_n_650));
  ON21X1 add_463_14_g1013(.A (add_463_14_n_662), .B (add_463_14_n_891),
       .C (add_463_14_n_896), .Q (add_463_14_n_653));
  INX1 add_463_14_g1014(.A (add_463_14_n_654), .Q (add_463_14_n_655));
  EN2X0 add_463_14_g1016(.A (add_463_14_n_662), .B (add_463_14_n_814),
       .Q (n_6168));
  EN2X0 add_463_14_g1017(.A (add_463_14_n_664), .B (add_463_14_n_782),
       .Q (n_6170));
  EN2X0 add_463_14_g1018(.A (add_463_14_n_667), .B (add_463_14_n_808),
       .Q (n_6172));
  EN2X1 add_463_14_g1019(.A (add_463_14_n_669), .B (add_463_14_n_824),
       .Q (n_6174));
  INX1 add_463_14_g1020(.A (add_463_14_n_662), .Q (add_463_14_n_663));
  AN21X1 add_463_14_g1021(.A (add_463_14_n_676), .B (add_463_14_n_760),
       .C (add_463_14_n_702), .Q (add_463_14_n_662));
  AN221X1 add_463_14_g1022(.A (add_463_14_n_849), .B
       (add_463_14_n_741), .C (add_463_14_n_849), .D
       (add_463_14_n_676), .E (add_463_14_n_902), .Q
       (add_463_14_n_664));
  NO2X1 add_463_14_g1023(.A (add_463_14_n_676), .B (add_463_14_n_741),
       .Q (add_463_14_n_667));
  ON21X1 add_463_14_g1024(.A (n_6622), .B (add_463_14_n_889), .C
       (add_463_14_n_895), .Q (add_463_14_n_669));
  EN2X0 add_463_14_g1025(.A (add_463_14_n_679), .B (add_463_14_n_819),
       .Q (n_6178));
  EN2X0 add_463_14_g1026(.A (n_6622), .B (add_463_14_n_811), .Q
       (n_6176));
  AO221X1 add_463_14_g1027(.A (add_463_14_n_724), .B
       (add_463_14_n_695), .C (add_463_14_n_856), .D
       (add_463_14_n_739), .E (add_463_14_n_836), .Q
       (add_463_14_n_673));
  NO3X1 add_463_14_g1028(.A (n_6622), .B (add_463_14_n_889), .C
       (add_463_14_n_897), .Q (add_463_14_n_676));
  EN2X1 add_463_14_g1029(.A (add_463_14_n_696), .B (add_463_14_n_810),
       .Q (n_6180));
  AN21X1 add_463_14_g1030(.A (add_463_14_n_696), .B (add_463_14_n_890),
       .C (add_463_14_n_893), .Q (add_463_14_n_679));
  ON221X1 add_463_14_g1032(.A (add_463_14_n_722), .B
       (add_463_14_n_698), .C (add_463_14_n_888), .D
       (add_463_14_n_738), .E (add_463_14_n_885), .Q
       (add_463_14_n_683));
  OA21X1 add_463_14_g1033(.A (add_463_14_n_698), .B (add_463_14_n_762),
       .C (add_463_14_n_738), .Q (add_463_14_n_685));
  ON21X1 add_463_14_g1034(.A (add_463_14_n_698), .B (add_463_14_n_858),
       .C (add_463_14_n_839), .Q (add_463_14_n_687));
  AO221X1 add_463_14_g1035(.A (add_463_14_n_723), .B
       (add_463_14_n_705), .C (add_463_14_n_850), .D
       (add_463_14_n_744), .E (add_463_14_n_835), .Q
       (add_463_14_n_688));
  AO221X1 add_463_14_g1036(.A (add_463_14_n_719), .B
       (add_463_14_n_708), .C (add_463_14_n_857), .D
       (add_463_14_n_740), .E (add_463_14_n_844), .Q
       (add_463_14_n_691));
  INX1 add_463_14_g1037(.A (add_463_14_n_694), .Q (add_463_14_n_695));
  AN221X1 add_463_14_g1038(.A (add_463_14_n_761), .B
       (add_463_14_n_744), .C (add_463_14_n_721), .D
       (add_463_14_n_705), .E (add_463_14_n_748), .Q
       (add_463_14_n_694));
  FAX1 add_463_14_g1039(.A (n_6716), .B (n_6629), .CI
       (add_463_14_n_937), .S (n_6182), .CO (add_463_14_n_696));
  AN221X1 add_463_14_g1040(.A (add_463_14_n_836), .B
       (add_463_14_n_840), .C (add_463_14_n_756), .D
       (add_463_14_n_739), .E (add_463_14_n_833), .Q
       (add_463_14_n_698));
  AO221X1 add_463_14_g1041(.A (add_463_14_n_757), .B
       (add_463_14_n_740), .C (add_463_14_n_844), .D
       (add_463_14_n_845), .E (add_463_14_n_830), .Q
       (add_463_14_n_700));
  AO221X1 add_463_14_g1042(.A (add_463_14_n_741), .B
       (add_463_14_n_760), .C (add_463_14_n_902), .D
       (add_463_14_n_842), .E (add_463_14_n_878), .Q
       (add_463_14_n_702));
  INX1 add_463_14_g1043(.A (add_463_14_n_706), .Q (add_463_14_n_705));
  AN221X1 add_463_14_g1044(.A (add_463_14_n_901), .B
       (add_463_14_n_848), .C (add_463_14_n_742), .D
       (add_463_14_n_759), .E (add_463_14_n_832), .Q
       (add_463_14_n_706));
  AO221X1 add_463_14_g1045(.A (add_463_14_n_743), .B
       (add_463_14_n_758), .C (add_463_14_n_847), .D
       (add_463_14_n_904), .E (add_463_14_n_883), .Q
       (add_463_14_n_708));
  NO2X1 add_463_14_g1046(.A (add_463_14_n_727), .B (add_463_14_n_722),
       .Q (add_463_14_n_710));
  OR2X1 add_463_14_g1047(.A (add_463_14_n_727), .B (add_463_14_n_762),
       .Q (add_463_14_n_712));
  NO2X1 add_463_14_g1048(.A (add_463_14_n_727), .B (add_463_14_n_858),
       .Q (add_463_14_n_714));
  INX1 add_463_14_g1049(.A (add_463_14_n_716), .Q (add_463_14_n_717));
  NA2X1 add_463_14_g1050(.A (add_463_14_n_721), .B (add_463_14_n_725),
       .Q (add_463_14_n_716));
  INX1 add_463_14_g1051(.A (add_463_14_n_725), .Q (add_463_14_n_726));
  AND2X1 add_463_14_g1052(.A (add_463_14_n_765), .B (add_463_14_n_857),
       .Q (add_463_14_n_719));
  AND2X1 add_463_14_g1053(.A (add_463_14_n_757), .B (add_463_14_n_765),
       .Q (add_463_14_n_720));
  AND2X1 add_463_14_g1054(.A (add_463_14_n_761), .B (add_463_14_n_763),
       .Q (add_463_14_n_721));
  OR2X1 add_463_14_g1055(.A (add_463_14_n_762), .B (add_463_14_n_888),
       .Q (add_463_14_n_722));
  AND2X1 add_463_14_g1056(.A (add_463_14_n_763), .B (add_463_14_n_850),
       .Q (add_463_14_n_723));
  AND2X1 add_463_14_g1057(.A (add_463_14_n_764), .B (add_463_14_n_856),
       .Q (add_463_14_n_724));
  AND2X1 add_463_14_g1058(.A (add_463_14_n_759), .B (add_463_14_n_796),
       .Q (add_463_14_n_725));
  NA2X1 add_463_14_g1059(.A (add_463_14_n_756), .B (add_463_14_n_764),
       .Q (add_463_14_n_727));
  AND2X1 add_463_14_g1060(.A (add_463_14_n_758), .B (add_463_14_n_795),
       .Q (add_463_14_n_728));
  ON21X1 add_463_14_g1062(.A (add_463_14_n_838), .B (add_463_14_n_834),
       .C (add_463_14_n_829), .Q (add_463_14_n_748));
  OA21X1 add_463_14_g1063(.A (add_463_14_n_837), .B (add_463_14_n_839),
       .C (add_463_14_n_831), .Q (add_463_14_n_738));
  ON21X1 add_463_14_g1064(.A (add_463_14_n_843), .B (add_463_14_n_903),
       .C (add_463_14_n_884), .Q (add_463_14_n_739));
  ON21X1 add_463_14_g1065(.A (add_463_14_n_846), .B (add_463_14_n_905),
       .C (add_463_14_n_880), .Q (add_463_14_n_740));
  ON21X1 add_463_14_g1066(.A (add_463_14_n_895), .B (add_463_14_n_897),
       .C (add_463_14_n_877), .Q (add_463_14_n_741));
  ON21X1 add_463_14_g1067(.A (add_463_14_n_894), .B (add_463_14_n_898),
       .C (add_463_14_n_881), .Q (add_463_14_n_742));
  ON21X1 add_463_14_g1068(.A (add_463_14_n_896), .B (add_463_14_n_899),
       .C (add_463_14_n_879), .Q (add_463_14_n_743));
  ON21X1 add_463_14_g1069(.A (add_463_14_n_841), .B (add_463_14_n_887),
       .C (add_463_14_n_886), .Q (add_463_14_n_744));
  NA2I1X1 add_463_14_g1070(.B (add_463_14_n_847), .AN
       (add_463_14_n_883), .Q (add_463_14_n_766));
  AND2X1 add_463_14_g1071(.A (add_463_14_n_840), .B (add_463_14_n_856),
       .Q (add_463_14_n_756));
  AND2X1 add_463_14_g1072(.A (add_463_14_n_845), .B (add_463_14_n_857),
       .Q (add_463_14_n_757));
  NO2I1X1 add_463_14_g1073(.B (add_463_14_n_838), .AN
       (add_463_14_n_829), .Q (add_463_14_n_771));
  NO2I1X1 add_463_14_g1074(.B (add_463_14_n_830), .AN
       (add_463_14_n_845), .Q (add_463_14_n_774));
  NO2I1X1 add_463_14_g1075(.B (add_463_14_n_833), .AN
       (add_463_14_n_840), .Q (add_463_14_n_776));
  AND2X1 add_463_14_g1076(.A (add_463_14_n_847), .B (add_463_14_n_853),
       .Q (add_463_14_n_758));
  AND2X1 add_463_14_g1077(.A (add_463_14_n_848), .B (add_463_14_n_855),
       .Q (add_463_14_n_759));
  AND2X1 add_463_14_g1078(.A (add_463_14_n_842), .B (add_463_14_n_849),
       .Q (add_463_14_n_760));
  NA2I1X1 add_463_14_g1079(.B (add_463_14_n_885), .AN
       (add_463_14_n_888), .Q (add_463_14_n_780));
  NO2I1X1 add_463_14_g1080(.B (add_463_14_n_838), .AN
       (add_463_14_n_850), .Q (add_463_14_n_761));
  NO2I1X1 add_463_14_g1081(.B (add_463_14_n_878), .AN
       (add_463_14_n_842), .Q (add_463_14_n_782));
  NA2I1X1 add_463_14_g1082(.B (add_463_14_n_839), .AN
       (add_463_14_n_858), .Q (add_463_14_n_784));
  NO2I1X1 add_463_14_g1083(.B (add_463_14_n_837), .AN
       (add_463_14_n_831), .Q (add_463_14_n_785));
  NO2I1X1 add_463_14_g1084(.B (add_463_14_n_836), .AN
       (add_463_14_n_856), .Q (add_463_14_n_788));
  AND2X1 add_463_14_g1085(.A (add_463_14_n_850), .B (add_463_14_n_834),
       .Q (add_463_14_n_789));
  NO2I1X1 add_463_14_g1086(.B (add_463_14_n_844), .AN
       (add_463_14_n_857), .Q (add_463_14_n_791));
  OR2X1 add_463_14_g1087(.A (add_463_14_n_858), .B (add_463_14_n_837),
       .Q (add_463_14_n_762));
  NO2X1 add_463_14_g1088(.A (add_463_14_n_851), .B (add_463_14_n_841),
       .Q (add_463_14_n_763));
  NO2X1 add_463_14_g1089(.A (add_463_14_n_854), .B (add_463_14_n_843),
       .Q (add_463_14_n_764));
  NO2I1X1 add_463_14_g1090(.B (add_463_14_n_846), .AN
       (add_463_14_n_852), .Q (add_463_14_n_765));
  EO2X1 add_463_14_g1091(.A (\rs1_data[0]_39306 ), .B (n_6014), .Q
       (n_6184));
  NA2X1 add_463_14_g1092(.A (add_463_14_n_852), .B (add_463_14_n_905),
       .Q (add_463_14_n_798));
  NA2I1X1 add_463_14_g1093(.B (add_463_14_n_886), .AN
       (add_463_14_n_841), .Q (add_463_14_n_800));
  NO2I1X1 add_463_14_g1094(.B (add_463_14_n_851), .AN
       (add_463_14_n_887), .Q (add_463_14_n_802));
  NA2I1X1 add_463_14_g1095(.B (add_463_14_n_880), .AN
       (add_463_14_n_846), .Q (add_463_14_n_803));
  NA2I1X1 add_463_14_g1096(.B (add_463_14_n_884), .AN
       (add_463_14_n_843), .Q (add_463_14_n_805));
  NO2I1X1 add_463_14_g1097(.B (add_463_14_n_901), .AN
       (add_463_14_n_855), .Q (add_463_14_n_807));
  NO2I1X1 add_463_14_g1098(.B (add_463_14_n_902), .AN
       (add_463_14_n_849), .Q (add_463_14_n_808));
  NO2I1X1 add_463_14_g1099(.B (add_463_14_n_854), .AN
       (add_463_14_n_903), .Q (add_463_14_n_809));
  NA2I1X1 add_463_14_g1100(.B (add_463_14_n_890), .AN
       (add_463_14_n_893), .Q (add_463_14_n_810));
  NO2I1X1 add_463_14_g1101(.B (add_463_14_n_889), .AN
       (add_463_14_n_895), .Q (add_463_14_n_811));
  NA2I1X1 add_463_14_g1102(.B (add_463_14_n_894), .AN
       (add_463_14_n_892), .Q (add_463_14_n_812));
  NO2I1X1 add_463_14_g1103(.B (add_463_14_n_891), .AN
       (add_463_14_n_896), .Q (add_463_14_n_814));
  NO2I1X1 add_463_14_g1104(.B (add_463_14_n_904), .AN
       (add_463_14_n_853), .Q (add_463_14_n_816));
  NO2I1X1 add_463_14_g1105(.B (add_463_14_n_832), .AN
       (add_463_14_n_848), .Q (add_463_14_n_817));
  NO2I1X1 add_463_14_g1106(.B (add_463_14_n_882), .AN
       (add_463_14_n_900), .Q (add_463_14_n_819));
  NA2I1X1 add_463_14_g1107(.B (add_463_14_n_881), .AN
       (add_463_14_n_898), .Q (add_463_14_n_821));
  NA2I1X1 add_463_14_g1108(.B (add_463_14_n_877), .AN
       (add_463_14_n_897), .Q (add_463_14_n_824));
  NA2I1X1 add_463_14_g1109(.B (add_463_14_n_879), .AN
       (add_463_14_n_899), .Q (add_463_14_n_826));
  NO2X1 add_463_14_g1110(.A (add_463_14_n_891), .B (add_463_14_n_899),
       .Q (add_463_14_n_795));
  NO2X1 add_463_14_g1111(.A (add_463_14_n_892), .B (add_463_14_n_898),
       .Q (add_463_14_n_796));
  INX1 add_463_14_g1112(.A (add_463_14_n_834), .Q (add_463_14_n_835));
  NA2X1 add_463_14_g1113(.A (\rs1_data[23]_39246 ), .B (n_6000), .Q
       (add_463_14_n_829));
  AND2X1 add_463_14_g1114(.A (\rs1_data[15]_39476 ), .B (n_6005), .Q
       (add_463_14_n_830));
  NA2X1 add_463_14_g1115(.A (\rs1_data[29]_39336 ), .B (n_5994), .Q
       (add_463_14_n_831));
  AND2X1 add_463_14_g1116(.A (n_4477), .B (n_6001), .Q
       (add_463_14_n_832));
  AND2X1 add_463_14_g1117(.A (\rs1_data[27]_39286 ), .B (n_5996), .Q
       (add_463_14_n_833));
  NA2X1 add_463_14_g1118(.A (n_4463), .B (n_5991), .Q
       (add_463_14_n_834));
  AND2X1 add_463_14_g1119(.A (\rs1_data[26]_39276 ), .B (n_5997), .Q
       (add_463_14_n_836));
  NO2X1 add_463_14_g1120(.A (\rs1_data[29]_39336 ), .B (n_5994), .Q
       (add_463_14_n_837));
  NO2X1 add_463_14_g1121(.A (\rs1_data[23]_39246 ), .B (n_6000), .Q
       (add_463_14_n_838));
  NA2X1 add_463_14_g1122(.A (\rs1_data[28]_39296 ), .B (n_5995), .Q
       (add_463_14_n_839));
  OR2X1 add_463_14_g1123(.A (\rs1_data[27]_39286 ), .B (n_5996), .Q
       (add_463_14_n_840));
  NO2X1 add_463_14_g1124(.A (n_4479), .B (n_6015), .Q
       (add_463_14_n_841));
  OR2X1 add_463_14_g1125(.A (n_4460), .B (n_6556), .Q
       (add_463_14_n_842));
  NO2X1 add_463_14_g1126(.A (n_4481), .B (n_5998), .Q
       (add_463_14_n_843));
  AND2X1 add_463_14_g1127(.A (\rs1_data[14]_39466 ), .B (n_6006), .Q
       (add_463_14_n_844));
  OR2X1 add_463_14_g1128(.A (\rs1_data[15]_39476 ), .B (n_6005), .Q
       (add_463_14_n_845));
  NO2X1 add_463_14_g1129(.A (n_4476), .B (n_6007), .Q
       (add_463_14_n_846));
  OR2X1 add_463_14_g1130(.A (n_4474), .B (n_6013), .Q
       (add_463_14_n_847));
  OR2X1 add_463_14_g1131(.A (n_4477), .B (n_6001), .Q
       (add_463_14_n_848));
  OR2X1 add_463_14_g1132(.A (n_4466), .B (n_6555), .Q
       (add_463_14_n_849));
  OR2X1 add_463_14_g1133(.A (n_4463), .B (n_5991), .Q
       (add_463_14_n_850));
  NO2X1 add_463_14_g1134(.A (n_4486), .B (n_5992), .Q
       (add_463_14_n_851));
  OR2X1 add_463_14_g1135(.A (n_4475), .B (n_6008), .Q
       (add_463_14_n_852));
  OR2X1 add_463_14_g1136(.A (n_4480), .B (n_6559), .Q
       (add_463_14_n_853));
  NO2X1 add_463_14_g1137(.A (n_4483), .B (n_5999), .Q
       (add_463_14_n_854));
  OR2X1 add_463_14_g1138(.A (n_4478), .B (n_6002), .Q
       (add_463_14_n_855));
  OR2X1 add_463_14_g1139(.A (\rs1_data[26]_39276 ), .B (n_5997), .Q
       (add_463_14_n_856));
  OR2X1 add_463_14_g1140(.A (\rs1_data[14]_39466 ), .B (n_6006), .Q
       (add_463_14_n_857));
  NO2X1 add_463_14_g1141(.A (\rs1_data[28]_39296 ), .B (n_5995), .Q
       (add_463_14_n_858));
  INX1 add_463_14_g1142(.A (add_463_14_n_905), .Q (add_463_14_n_906));
  NA2X1 add_463_14_g1143(.A (n_4461), .B (n_6554), .Q
       (add_463_14_n_877));
  AND2X1 add_463_14_g1144(.A (n_4460), .B (n_6556), .Q
       (add_463_14_n_878));
  NA2X1 add_463_14_g1145(.A (n_4487), .B (n_6558), .Q
       (add_463_14_n_879));
  NA2X1 add_463_14_g1146(.A (n_4476), .B (n_6007), .Q
       (add_463_14_n_880));
  NA2X1 add_463_14_g1147(.A (n_4482), .B (n_6003), .Q
       (add_463_14_n_881));
  AND2X1 add_463_14_g1148(.A (n_6757), .B (n_6010), .Q
       (add_463_14_n_882));
  AND2X1 add_463_14_g1149(.A (n_4474), .B (n_6013), .Q
       (add_463_14_n_883));
  NA2X1 add_463_14_g1150(.A (n_4481), .B (n_5998), .Q
       (add_463_14_n_884));
  NA2X1 add_463_14_g1151(.A (n_4485), .B (n_5993), .Q
       (add_463_14_n_885));
  NA2X1 add_463_14_g1152(.A (n_4479), .B (n_6015), .Q
       (add_463_14_n_886));
  NA2X1 add_463_14_g1153(.A (n_4486), .B (n_5992), .Q
       (add_463_14_n_887));
  NO2X1 add_463_14_g1154(.A (n_4485), .B (n_5993), .Q
       (add_463_14_n_888));
  NO2X1 add_463_14_g1155(.A (n_4465), .B (n_6717), .Q
       (add_463_14_n_889));
  OR2X1 add_463_14_g1156(.A (n_6628), .B (n_6011), .Q
       (add_463_14_n_890));
  NO2X1 add_463_14_g1157(.A (n_4464), .B (n_6557), .Q
       (add_463_14_n_891));
  NO2X1 add_463_14_g1158(.A (n_4484), .B (n_6004), .Q
       (add_463_14_n_892));
  AND2X1 add_463_14_g1159(.A (n_6628), .B (n_6011), .Q
       (add_463_14_n_893));
  NA2X1 add_463_14_g1160(.A (n_4484), .B (n_6004), .Q
       (add_463_14_n_894));
  NA2X1 add_463_14_g1161(.A (n_4465), .B (n_6717), .Q
       (add_463_14_n_895));
  NA2X1 add_463_14_g1162(.A (n_4464), .B (n_6557), .Q
       (add_463_14_n_896));
  NO2X1 add_463_14_g1163(.A (n_4461), .B (n_6554), .Q
       (add_463_14_n_897));
  NO2X1 add_463_14_g1164(.A (n_4482), .B (n_6003), .Q
       (add_463_14_n_898));
  NO2X1 add_463_14_g1165(.A (n_4487), .B (n_6558), .Q
       (add_463_14_n_899));
  OR2X1 add_463_14_g1166(.A (n_6757), .B (n_6010), .Q
       (add_463_14_n_900));
  AND2X1 add_463_14_g1168(.A (n_4478), .B (n_6002), .Q
       (add_463_14_n_901));
  AND2X1 add_463_14_g1169(.A (n_4466), .B (n_6555), .Q
       (add_463_14_n_902));
  NA2X1 add_463_14_g1170(.A (n_4483), .B (n_5999), .Q
       (add_463_14_n_903));
  AND2X1 add_463_14_g1171(.A (n_4480), .B (n_6559), .Q
       (add_463_14_n_904));
  NA2X1 add_463_14_g1172(.A (n_4475), .B (n_6008), .Q
       (add_463_14_n_905));
  AND2X1 add_463_14_g1174(.A (\rs1_data[0]_39306 ), .B (n_6014), .Q
       (add_463_14_n_937));
  EN3X1 add_463_14_g1176(.A (add_463_14_n_610), .B
       (alu_sra_result[31]), .C (n_6560), .Q (n_6122));
  AO321X1 add_463_14_g1178(.A (add_463_14_n_728), .B
       (add_463_14_n_720), .C (add_463_14_n_663), .D
       (add_463_14_n_720), .E (add_463_14_n_708), .F
       (add_463_14_n_700), .Q (add_463_14_n_654));
  MU2IX1 inc_ADD_UNS_OP_5_g2724(.S (inc_ADD_UNS_OP_5_n_2648), .IN0
       (csr_minstret[62]), .IN1 (inc_ADD_UNS_OP_5_n_2929), .Q (n_5756));
  NA2X1 inc_ADD_UNS_OP_5_g2727(.A (inc_ADD_UNS_OP_5_n_2656), .B
       (inc_ADD_UNS_OP_5_n_2889), .Q (inc_ADD_UNS_OP_5_n_2648));
  NA2X1 inc_ADD_UNS_OP_5_g2730(.A (inc_ADD_UNS_OP_5_n_2661), .B
       (inc_ADD_UNS_OP_5_n_2894), .Q (inc_ADD_UNS_OP_5_n_2652));
  MU2IX1 inc_ADD_UNS_OP_5_g2731(.S (inc_ADD_UNS_OP_5_n_2665), .IN0
       (csr_minstret[58]), .IN1 (inc_ADD_UNS_OP_5_n_2970), .Q (n_5760));
  NO2X1 inc_ADD_UNS_OP_5_g2733(.A (inc_ADD_UNS_OP_5_n_2665), .B
       (inc_ADD_UNS_OP_5_n_2970), .Q (inc_ADD_UNS_OP_5_n_2656));
  MU2IX1 inc_ADD_UNS_OP_5_g2734(.S (inc_ADD_UNS_OP_5_n_2667), .IN0
       (csr_minstret[60]), .IN1 (inc_ADD_UNS_OP_5_n_2966), .Q (n_5758));
  NO2X2 inc_ADD_UNS_OP_5_g2735(.A (inc_ADD_UNS_OP_5_n_2667), .B
       (inc_ADD_UNS_OP_5_n_2966), .Q (inc_ADD_UNS_OP_5_n_2661));
  NA2X2 inc_ADD_UNS_OP_5_g2737(.A (inc_ADD_UNS_OP_5_n_2672), .B
       (csr_minstret[57]), .Q (inc_ADD_UNS_OP_5_n_2665));
  NA2X2 inc_ADD_UNS_OP_5_g2738(.A (inc_ADD_UNS_OP_5_n_2672), .B
       (inc_ADD_UNS_OP_5_n_2886), .Q (inc_ADD_UNS_OP_5_n_2667));
  MU2IX1 inc_ADD_UNS_OP_5_g2740(.S (inc_ADD_UNS_OP_5_n_2678), .IN0
       (csr_minstret[56]), .IN1 (inc_ADD_UNS_OP_5_n_2931), .Q (n_5762));
  NO2X2 inc_ADD_UNS_OP_5_g2742(.A (inc_ADD_UNS_OP_5_n_2678), .B
       (inc_ADD_UNS_OP_5_n_2931), .Q (inc_ADD_UNS_OP_5_n_2672));
  NA2X2 inc_ADD_UNS_OP_5_g2744(.A (inc_ADD_UNS_OP_5_n_2683), .B
       (csr_minstret[55]), .Q (inc_ADD_UNS_OP_5_n_2678));
  AND6X2 inc_ADD_UNS_OP_5_g2748(.A (inc_ADD_UNS_OP_5_n_2710), .B
       (csr_minstret[50]), .C (csr_minstret[52]), .D
       (csr_minstret[51]), .E (csr_minstret[53]), .F
       (csr_minstret[54]), .Q (inc_ADD_UNS_OP_5_n_2683));
  NA2X1 inc_ADD_UNS_OP_5_g2750(.A (inc_ADD_UNS_OP_5_n_2693), .B
       (csr_minstret[53]), .Q (inc_ADD_UNS_OP_5_n_2688));
  MU2IX1 inc_ADD_UNS_OP_5_g2752(.S (inc_ADD_UNS_OP_5_n_2699), .IN0
       (csr_minstret[52]), .IN1 (inc_ADD_UNS_OP_5_n_2948), .Q (n_5766));
  NO2X1 inc_ADD_UNS_OP_5_g2753(.A (inc_ADD_UNS_OP_5_n_2699), .B
       (inc_ADD_UNS_OP_5_n_2948), .Q (inc_ADD_UNS_OP_5_n_2693));
  NA2X1 inc_ADD_UNS_OP_5_g2755(.A (inc_ADD_UNS_OP_5_n_2704), .B
       (csr_minstret[51]), .Q (inc_ADD_UNS_OP_5_n_2699));
  MU2IX1 inc_ADD_UNS_OP_5_g2757(.S (inc_ADD_UNS_OP_5_n_2708), .IN0
       (csr_minstret[50]), .IN1 (inc_ADD_UNS_OP_5_n_2924), .Q (n_5768));
  NO2X1 inc_ADD_UNS_OP_5_g2759(.A (inc_ADD_UNS_OP_5_n_2708), .B
       (inc_ADD_UNS_OP_5_n_2924), .Q (inc_ADD_UNS_OP_5_n_2704));
  INX1 inc_ADD_UNS_OP_5_g2761(.A (inc_ADD_UNS_OP_5_n_2710), .Q
       (inc_ADD_UNS_OP_5_n_2708));
  AND6X2 inc_ADD_UNS_OP_5_g2765(.A (inc_ADD_UNS_OP_5_n_2730), .B
       (csr_minstret[45]), .C (csr_minstret[47]), .D
       (csr_minstret[46]), .E (csr_minstret[48]), .F
       (csr_minstret[49]), .Q (inc_ADD_UNS_OP_5_n_2710));
  NA2X1 inc_ADD_UNS_OP_5_g2767(.A (inc_ADD_UNS_OP_5_n_2720), .B
       (csr_minstret[48]), .Q (inc_ADD_UNS_OP_5_n_2718));
  HAX2 inc_ADD_UNS_OP_5_g2769(.A (inc_ADD_UNS_OP_5_n_2724), .B
       (csr_minstret[47]), .S (n_5771), .CO (inc_ADD_UNS_OP_5_n_2720));
  HAX2 inc_ADD_UNS_OP_5_g2770(.A (inc_ADD_UNS_OP_5_n_2727), .B
       (csr_minstret[46]), .S (n_5772), .CO (inc_ADD_UNS_OP_5_n_2724));
  HAX2 inc_ADD_UNS_OP_5_g2771(.A (inc_ADD_UNS_OP_5_n_2730), .B
       (csr_minstret[45]), .S (n_5773), .CO (inc_ADD_UNS_OP_5_n_2727));
  AND6X2 inc_ADD_UNS_OP_5_g2775(.A (inc_ADD_UNS_OP_5_n_2752), .B
       (csr_minstret[40]), .C (csr_minstret[42]), .D
       (csr_minstret[41]), .E (csr_minstret[43]), .F
       (csr_minstret[44]), .Q (inc_ADD_UNS_OP_5_n_2730));
  NA2X1 inc_ADD_UNS_OP_5_g2777(.A (inc_ADD_UNS_OP_5_n_2740), .B
       (csr_minstret[43]), .Q (inc_ADD_UNS_OP_5_n_2738));
  HAX2 inc_ADD_UNS_OP_5_g2779(.A (inc_ADD_UNS_OP_5_n_2744), .B
       (csr_minstret[42]), .S (n_5776), .CO (inc_ADD_UNS_OP_5_n_2740));
  HAX2 inc_ADD_UNS_OP_5_g2780(.A (inc_ADD_UNS_OP_5_n_2747), .B
       (csr_minstret[41]), .S (n_5777), .CO (inc_ADD_UNS_OP_5_n_2744));
  HAX2 inc_ADD_UNS_OP_5_g2781(.A (inc_ADD_UNS_OP_5_n_2752), .B
       (csr_minstret[40]), .S (n_5778), .CO (inc_ADD_UNS_OP_5_n_2747));
  AND6X2 inc_ADD_UNS_OP_5_g2783(.A (inc_ADD_UNS_OP_5_n_2770), .B
       (csr_minstret[35]), .C (csr_minstret[37]), .D
       (csr_minstret[36]), .E (csr_minstret[38]), .F
       (csr_minstret[39]), .Q (inc_ADD_UNS_OP_5_n_2752));
  NA2X1 inc_ADD_UNS_OP_5_g2785(.A (inc_ADD_UNS_OP_5_n_2758), .B
       (csr_minstret[38]), .Q (inc_ADD_UNS_OP_5_n_2756));
  HAX2 inc_ADD_UNS_OP_5_g2787(.A (inc_ADD_UNS_OP_5_n_2762), .B
       (csr_minstret[37]), .S (n_5781), .CO (inc_ADD_UNS_OP_5_n_2758));
  HAX2 inc_ADD_UNS_OP_5_g2788(.A (inc_ADD_UNS_OP_5_n_2765), .B
       (csr_minstret[36]), .S (n_5782), .CO (inc_ADD_UNS_OP_5_n_2762));
  HAX2 inc_ADD_UNS_OP_5_g2789(.A (inc_ADD_UNS_OP_5_n_2770), .B
       (csr_minstret[35]), .S (n_5783), .CO (inc_ADD_UNS_OP_5_n_2765));
  AND6X2 inc_ADD_UNS_OP_5_g2791(.A (inc_ADD_UNS_OP_5_n_2788), .B
       (n_5985), .C (n_5729), .D (csr_minstret[32]), .E
       (csr_minstret[33]), .F (csr_minstret[34]), .Q
       (inc_ADD_UNS_OP_5_n_2770));
  NA2X1 inc_ADD_UNS_OP_5_g2793(.A (inc_ADD_UNS_OP_5_n_2776), .B
       (csr_minstret[33]), .Q (inc_ADD_UNS_OP_5_n_2774));
  HAX1 inc_ADD_UNS_OP_5_g2795(.A (inc_ADD_UNS_OP_5_n_2780), .B
       (csr_minstret[32]), .S (n_5786), .CO (inc_ADD_UNS_OP_5_n_2776));
  HAX1 inc_ADD_UNS_OP_5_g2796(.A (inc_ADD_UNS_OP_5_n_2783), .B
       (n_5985), .S (n_5787), .CO (inc_ADD_UNS_OP_5_n_2780));
  HAX1 inc_ADD_UNS_OP_5_g2797(.A (inc_ADD_UNS_OP_5_n_2788), .B
       (n_5729), .S (n_5788), .CO (inc_ADD_UNS_OP_5_n_2783));
  EO2X1 inc_ADD_UNS_OP_5_g2798(.A (inc_ADD_UNS_OP_5_n_2791), .B
       (n_5730), .Q (n_5789));
  AND6X2 inc_ADD_UNS_OP_5_g2799(.A (inc_ADD_UNS_OP_5_n_2805), .B
       (n_5733), .C (n_5732), .D (n_5734), .E (n_5731), .F (n_5730), .Q
       (inc_ADD_UNS_OP_5_n_2788));
  HAX1 inc_ADD_UNS_OP_5_g2800(.A (inc_ADD_UNS_OP_5_n_2794), .B
       (n_5731), .S (n_5790), .CO (inc_ADD_UNS_OP_5_n_2791));
  HAX1 inc_ADD_UNS_OP_5_g2801(.A (inc_ADD_UNS_OP_5_n_2797), .B
       (n_5732), .S (n_5791), .CO (inc_ADD_UNS_OP_5_n_2794));
  HAX1 inc_ADD_UNS_OP_5_g2802(.A (inc_ADD_UNS_OP_5_n_2800), .B
       (n_5733), .S (n_5792), .CO (inc_ADD_UNS_OP_5_n_2797));
  HAX1 inc_ADD_UNS_OP_5_g2803(.A (inc_ADD_UNS_OP_5_n_2805), .B
       (n_5734), .S (n_5793), .CO (inc_ADD_UNS_OP_5_n_2800));
  EO2X1 inc_ADD_UNS_OP_5_g2804(.A (inc_ADD_UNS_OP_5_n_2808), .B
       (n_5735), .Q (n_5794));
  AND6X2 inc_ADD_UNS_OP_5_g2805(.A (inc_ADD_UNS_OP_5_n_2820), .B
       (n_5737), .C (n_5736), .D (n_5739), .E (n_5738), .F (n_5735), .Q
       (inc_ADD_UNS_OP_5_n_2805));
  HAX1 inc_ADD_UNS_OP_5_g2806(.A (inc_ADD_UNS_OP_5_n_2811), .B
       (n_5736), .S (n_5795), .CO (inc_ADD_UNS_OP_5_n_2808));
  HAX1 inc_ADD_UNS_OP_5_g2807(.A (inc_ADD_UNS_OP_5_n_2814), .B
       (n_5737), .S (n_5796), .CO (inc_ADD_UNS_OP_5_n_2811));
  HAX1 inc_ADD_UNS_OP_5_g2808(.A (inc_ADD_UNS_OP_5_n_2817), .B
       (n_5738), .S (n_5797), .CO (inc_ADD_UNS_OP_5_n_2814));
  HAX1 inc_ADD_UNS_OP_5_g2809(.A (inc_ADD_UNS_OP_5_n_2820), .B
       (n_5739), .S (n_5798), .CO (inc_ADD_UNS_OP_5_n_2817));
  HAX2 inc_ADD_UNS_OP_5_g2810(.A (inc_ADD_UNS_OP_5_n_2823), .B
       (n_5740), .S (n_5799), .CO (inc_ADD_UNS_OP_5_n_2820));
  HAX2 inc_ADD_UNS_OP_5_g2811(.A (inc_ADD_UNS_OP_5_n_2825), .B
       (n_5741), .S (n_5800), .CO (inc_ADD_UNS_OP_5_n_2823));
  EO2X1 inc_ADD_UNS_OP_5_g2812(.A (inc_ADD_UNS_OP_5_n_2828), .B
       (n_5742), .Q (n_5801));
  AND5X1 inc_ADD_UNS_OP_5_g2813(.A (inc_ADD_UNS_OP_5_n_2837), .B
       (n_4536), .C (n_4538), .D (n_5743), .E (n_5742), .Q
       (inc_ADD_UNS_OP_5_n_2825));
  HAX1 inc_ADD_UNS_OP_5_g2814(.A (inc_ADD_UNS_OP_5_n_2831), .B
       (n_5743), .S (n_5802), .CO (inc_ADD_UNS_OP_5_n_2828));
  HAX1 inc_ADD_UNS_OP_5_g2815(.A (inc_ADD_UNS_OP_5_n_2834), .B
       (n_4538), .S (n_5803), .CO (inc_ADD_UNS_OP_5_n_2831));
  HAX1 inc_ADD_UNS_OP_5_g2816(.A (inc_ADD_UNS_OP_5_n_2837), .B
       (n_4536), .S (n_5804), .CO (inc_ADD_UNS_OP_5_n_2834));
  HAX1 inc_ADD_UNS_OP_5_g2817(.A (inc_ADD_UNS_OP_5_n_2840), .B
       (n_5746), .S (n_5805), .CO (inc_ADD_UNS_OP_5_n_2837));
  HAX1 inc_ADD_UNS_OP_5_g2818(.A (inc_ADD_UNS_OP_5_n_2842), .B
       (n_5747), .S (n_5806), .CO (inc_ADD_UNS_OP_5_n_2840));
  HAX1 inc_ADD_UNS_OP_5_g2819(.A (inc_ADD_UNS_OP_5_n_2844), .B
       (n_5748), .S (n_5807), .CO (inc_ADD_UNS_OP_5_n_2842));
  EO2X1 inc_ADD_UNS_OP_5_g2820(.A (inc_ADD_UNS_OP_5_n_2847), .B
       (n_5749), .Q (n_5808));
  AND2X2 inc_ADD_UNS_OP_5_g2821(.A (inc_ADD_UNS_OP_5_n_2847), .B
       (n_5749), .Q (inc_ADD_UNS_OP_5_n_2844));
  HAX2 inc_ADD_UNS_OP_5_g2822(.A (inc_ADD_UNS_OP_5_n_2850), .B
       (n_5750), .S (n_5809), .CO (inc_ADD_UNS_OP_5_n_2847));
  EO2X1 inc_ADD_UNS_OP_5_g2823(.A (inc_ADD_UNS_OP_5_n_2855), .B
       (n_5751), .Q (n_5810));
  NO2I1X2 inc_ADD_UNS_OP_5_g2826(.B (inc_ADD_UNS_OP_5_n_2860), .AN
       (n_6726), .Q (inc_ADD_UNS_OP_5_n_2855));
  EO2X1 inc_ADD_UNS_OP_5_g2828(.A (inc_ADD_UNS_OP_5_n_2987), .B
       (n_6730), .Q (n_5812));
  NA2X1 inc_ADD_UNS_OP_5_g2829(.A (inc_ADD_UNS_OP_5_n_2987), .B
       (n_6730), .Q (inc_ADD_UNS_OP_5_n_2860));
  EO2X1 inc_ADD_UNS_OP_5_g2830(.A (inc_ADD_UNS_OP_5_n_2868), .B
       (n_6731), .Q (n_5813));
  HAX2 inc_ADD_UNS_OP_5_g2833(.A (inc_ADD_UNS_OP_5_n_2871), .B
       (n_4535), .S (n_5814), .CO (inc_ADD_UNS_OP_5_n_2868));
  EO2X1 inc_ADD_UNS_OP_5_g2837(.A (inc_ADD_UNS_OP_5_n_2881), .B
       (n_5988), .Q (n_5816));
  NA2X2 inc_ADD_UNS_OP_5_g2838(.A (inc_ADD_UNS_OP_5_n_2881), .B
       (n_5988), .Q (inc_ADD_UNS_OP_5_n_2876));
  NO2I1X1 inc_ADD_UNS_OP_5_g2840(.B (inc_ADD_UNS_OP_5_n_2891), .AN
       (n_6724), .Q (inc_ADD_UNS_OP_5_n_2881));
  EO2X1 inc_ADD_UNS_OP_5_g2842(.A (n_4534), .B (n_6239), .Q (n_5818));
  NO3X1 inc_ADD_UNS_OP_5_g2843(.A (inc_ADD_UNS_OP_5_n_2973), .B
       (inc_ADD_UNS_OP_5_n_2968), .C (inc_ADD_UNS_OP_5_n_2970), .Q
       (inc_ADD_UNS_OP_5_n_2886));
  NO3X1 inc_ADD_UNS_OP_5_g2844(.A (inc_ADD_UNS_OP_5_n_2966), .B
       (inc_ADD_UNS_OP_5_n_2974), .C (inc_ADD_UNS_OP_5_n_2968), .Q
       (inc_ADD_UNS_OP_5_n_2889));
  NA2X1 inc_ADD_UNS_OP_5_g2845(.A (n_4534), .B (n_6239), .Q
       (inc_ADD_UNS_OP_5_n_2891));
  NO2X1 inc_ADD_UNS_OP_5_g2846(.A (inc_ADD_UNS_OP_5_n_2974), .B
       (inc_ADD_UNS_OP_5_n_2929), .Q (inc_ADD_UNS_OP_5_n_2894));
  INX1 inc_ADD_UNS_OP_5_g2848(.A (csr_minstret[50]), .Q
       (inc_ADD_UNS_OP_5_n_2924));
  INX1 inc_ADD_UNS_OP_5_g2850(.A (csr_minstret[62]), .Q
       (inc_ADD_UNS_OP_5_n_2929));
  INX1 inc_ADD_UNS_OP_5_g2851(.A (csr_minstret[56]), .Q
       (inc_ADD_UNS_OP_5_n_2931));
  INX1 inc_ADD_UNS_OP_5_g2856(.A (csr_minstret[52]), .Q
       (inc_ADD_UNS_OP_5_n_2948));
  INX1 inc_ADD_UNS_OP_5_g2864(.A (csr_minstret[60]), .Q
       (inc_ADD_UNS_OP_5_n_2966));
  INX1 inc_ADD_UNS_OP_5_g2865(.A (csr_minstret[59]), .Q
       (inc_ADD_UNS_OP_5_n_2968));
  INX1 inc_ADD_UNS_OP_5_g2866(.A (csr_minstret[58]), .Q
       (inc_ADD_UNS_OP_5_n_2970));
  INX1 inc_ADD_UNS_OP_5_g2867(.A (csr_minstret[57]), .Q
       (inc_ADD_UNS_OP_5_n_2973));
  INX1 inc_ADD_UNS_OP_5_g2868(.A (csr_minstret[61]), .Q
       (inc_ADD_UNS_OP_5_n_2974));
  MU2IX1 inc_ADD_UNS_OP_5_g2(.S (inc_ADD_UNS_OP_5_n_2656), .IN0
       (inc_ADD_UNS_OP_5_n_2968), .IN1 (csr_minstret[59]), .Q (n_5759));
  MU2IX1 inc_ADD_UNS_OP_5_g2869(.S (inc_ADD_UNS_OP_5_n_2661), .IN0
       (inc_ADD_UNS_OP_5_n_2974), .IN1 (csr_minstret[61]), .Q (n_5757));
  MU2IX1 inc_ADD_UNS_OP_5_g2870(.S (inc_ADD_UNS_OP_5_n_2672), .IN0
       (inc_ADD_UNS_OP_5_n_2973), .IN1 (csr_minstret[57]), .Q (n_5761));
  EO2X1 inc_ADD_UNS_OP_5_g2871(.A (inc_ADD_UNS_OP_5_n_2683), .B
       (csr_minstret[55]), .Q (n_5763));
  EO2X1 inc_ADD_UNS_OP_5_g2872(.A (inc_ADD_UNS_OP_5_n_2693), .B
       (csr_minstret[53]), .Q (n_5765));
  EO2X1 inc_ADD_UNS_OP_5_g2873(.A (inc_ADD_UNS_OP_5_n_2704), .B
       (csr_minstret[51]), .Q (n_5767));
  EO2X1 inc_ADD_UNS_OP_5_g2874(.A (inc_ADD_UNS_OP_5_n_2720), .B
       (csr_minstret[48]), .Q (n_5770));
  EO2X1 inc_ADD_UNS_OP_5_g2875(.A (inc_ADD_UNS_OP_5_n_2740), .B
       (csr_minstret[43]), .Q (n_5775));
  EO2X1 inc_ADD_UNS_OP_5_g2876(.A (inc_ADD_UNS_OP_5_n_2758), .B
       (csr_minstret[38]), .Q (n_5780));
  EO2X1 inc_ADD_UNS_OP_5_g2877(.A (inc_ADD_UNS_OP_5_n_2776), .B
       (csr_minstret[33]), .Q (n_5785));
  EN2X1 inc_ADD_UNS_OP_5_g2878(.A (inc_ADD_UNS_OP_5_n_2860), .B
       (n_6726), .Q (n_5811));
  AND2X1 inc_ADD_UNS_OP_5_g2879(.A (inc_ADD_UNS_OP_5_n_2868), .B
       (n_6731), .Q (inc_ADD_UNS_OP_5_n_2987));
  EN2X1 inc_ADD_UNS_OP_5_g2880(.A (inc_ADD_UNS_OP_5_n_2876), .B
       (n_5987), .Q (n_5815));
  EN2X1 inc_ADD_UNS_OP_5_g2881(.A (inc_ADD_UNS_OP_5_n_2891), .B
       (n_6724), .Q (n_5817));
  EN2X1 inc_ADD_UNS_OP_5_g2882(.A (inc_ADD_UNS_OP_5_n_2652), .B
       (csr_minstret[63]), .Q (n_5755));
  EN2X1 inc_ADD_UNS_OP_5_g2883(.A (inc_ADD_UNS_OP_5_n_2688), .B
       (csr_minstret[54]), .Q (n_5764));
  EN2X1 inc_ADD_UNS_OP_5_g2884(.A (inc_ADD_UNS_OP_5_n_2718), .B
       (csr_minstret[49]), .Q (n_5769));
  EN2X1 inc_ADD_UNS_OP_5_g2885(.A (inc_ADD_UNS_OP_5_n_2756), .B
       (csr_minstret[39]), .Q (n_5779));
  EN2X1 inc_ADD_UNS_OP_5_g2886(.A (inc_ADD_UNS_OP_5_n_2774), .B
       (csr_minstret[34]), .Q (n_5784));
  EN2X1 inc_ADD_UNS_OP_5_g2887(.A (inc_ADD_UNS_OP_5_n_2738), .B
       (csr_minstret[44]), .Q (n_5774));
  AND2X2 inc_ADD_UNS_OP_5_g2889(.A (inc_ADD_UNS_OP_5_n_2855), .B
       (n_5751), .Q (inc_ADD_UNS_OP_5_n_2850));
  NO2I1X2 inc_ADD_UNS_OP_5_g2891(.B (inc_ADD_UNS_OP_5_n_2876), .AN
       (n_5987), .Q (inc_ADD_UNS_OP_5_n_2871));
  NA2X2 inc_add_1345_58_1_g819(.A (inc_add_1345_58_1_n_451), .B
       (n_5729), .Q (inc_add_1345_58_1_n_448));
  HAX2 inc_add_1345_58_1_g820(.A (inc_add_1345_58_1_n_454), .B
       (n_5730), .S (n_6308), .CO (inc_add_1345_58_1_n_451));
  HAX2 inc_add_1345_58_1_g821(.A (inc_add_1345_58_1_n_456), .B
       (n_5731), .S (n_6310), .CO (inc_add_1345_58_1_n_454));
  HAX2 inc_add_1345_58_1_g822(.A (inc_add_1345_58_1_n_458), .B
       (n_5732), .S (n_6312), .CO (inc_add_1345_58_1_n_456));
  HAX2 inc_add_1345_58_1_g823(.A (inc_add_1345_58_1_n_460), .B
       (n_5733), .S (n_6314), .CO (inc_add_1345_58_1_n_458));
  HAX2 inc_add_1345_58_1_g824(.A (inc_add_1345_58_1_n_462), .B
       (n_5734), .S (n_6316), .CO (inc_add_1345_58_1_n_460));
  HAX2 inc_add_1345_58_1_g825(.A (inc_add_1345_58_1_n_464), .B
       (n_5735), .S (n_6318), .CO (inc_add_1345_58_1_n_462));
  HAX2 inc_add_1345_58_1_g826(.A (inc_add_1345_58_1_n_466), .B
       (n_5736), .S (n_6320), .CO (inc_add_1345_58_1_n_464));
  NO2I1X4 inc_add_1345_58_1_g828(.B (inc_add_1345_58_1_n_471), .AN
       (n_5737), .Q (inc_add_1345_58_1_n_466));
  EO2X0 inc_add_1345_58_1_g830(.A (inc_add_1345_58_1_n_476), .B
       (n_5738), .Q (n_6335));
  NA2X1 inc_add_1345_58_1_g831(.A (inc_add_1345_58_1_n_476), .B
       (n_5738), .Q (inc_add_1345_58_1_n_471));
  NO2I1X4 inc_add_1345_58_1_g833(.B (inc_add_1345_58_1_n_481), .AN
       (n_5739), .Q (inc_add_1345_58_1_n_476));
  EO2X1 inc_add_1345_58_1_g835(.A (inc_add_1345_58_1_n_486), .B
       (n_5740), .Q (n_6350));
  NA2X1 inc_add_1345_58_1_g836(.A (inc_add_1345_58_1_n_486), .B
       (n_5740), .Q (inc_add_1345_58_1_n_481));
  EO2X0 inc_add_1345_58_1_g837(.A (inc_add_1345_58_1_n_728), .B
       (n_5741), .Q (n_6352));
  AND2X4 inc_add_1345_58_1_g838(.A (inc_add_1345_58_1_n_728), .B
       (n_5741), .Q (inc_add_1345_58_1_n_486));
  EO2X0 inc_add_1345_58_1_g839(.A (inc_add_1345_58_1_n_494), .B
       (n_5742), .Q (n_6354));
  HAX2 inc_add_1345_58_1_g842(.A (inc_add_1345_58_1_n_497), .B
       (n_5743), .S (n_6356), .CO (inc_add_1345_58_1_n_494));
  HAX2 inc_add_1345_58_1_g843(.A (inc_add_1345_58_1_n_499), .B
       (n_4538), .S (n_6358), .CO (inc_add_1345_58_1_n_497));
  NO2I1X4 inc_add_1345_58_1_g845(.B (inc_add_1345_58_1_n_504), .AN
       (n_4536), .Q (inc_add_1345_58_1_n_499));
  EO2X0 inc_add_1345_58_1_g847(.A (inc_add_1345_58_1_n_509), .B
       (n_5746), .Q (n_6362));
  NA2X2 inc_add_1345_58_1_g848(.A (inc_add_1345_58_1_n_509), .B
       (n_5746), .Q (inc_add_1345_58_1_n_504));
  EO2X0 inc_add_1345_58_1_g852(.A (inc_add_1345_58_1_n_517), .B
       (n_5748), .Q (n_6366));
  NA2X1 inc_add_1345_58_1_g853(.A (inc_add_1345_58_1_n_517), .B
       (n_5748), .Q (inc_add_1345_58_1_n_514));
  HAX2 inc_add_1345_58_1_g854(.A (inc_add_1345_58_1_n_520), .B
       (n_5749), .S (n_6369), .CO (inc_add_1345_58_1_n_517));
  EO2X1 inc_add_1345_58_1_g855(.A (inc_add_1345_58_1_n_525), .B
       (n_5750), .Q (n_6371));
  AND2X1 inc_add_1345_58_1_g856(.A (inc_add_1345_58_1_n_525), .B
       (n_5750), .Q (inc_add_1345_58_1_n_520));
  EO2X1 inc_add_1345_58_1_g857(.A (inc_add_1345_58_1_n_528), .B
       (n_5751), .Q (n_6374));
  AND4X1 inc_add_1345_58_1_g858(.A (inc_add_1345_58_1_n_534), .B
       (n_6730), .C (n_6726), .D (n_5751), .Q
       (inc_add_1345_58_1_n_525));
  HAX1 inc_add_1345_58_1_g859(.A (inc_add_1345_58_1_n_531), .B
       (n_6726), .S (n_6376), .CO (inc_add_1345_58_1_n_528));
  HAX1 inc_add_1345_58_1_g860(.A (inc_add_1345_58_1_n_534), .B
       (n_6730), .S (n_6378), .CO (inc_add_1345_58_1_n_531));
  HAX1 inc_add_1345_58_1_g861(.A (inc_add_1345_58_1_n_537), .B
       (n_6731), .S (n_6380), .CO (inc_add_1345_58_1_n_534));
  HAX1 inc_add_1345_58_1_g862(.A (inc_add_1345_58_1_n_539), .B
       (n_4535), .S (n_6382), .CO (inc_add_1345_58_1_n_537));
  EO2X0 inc_add_1345_58_1_g863(.A (inc_add_1345_58_1_n_544), .B
       (n_5987), .Q (n_6384));
  AND2X2 inc_add_1345_58_1_g864(.A (inc_add_1345_58_1_n_544), .B
       (n_5987), .Q (inc_add_1345_58_1_n_539));
  EO2X1 inc_add_1345_58_1_g865(.A (inc_add_1345_58_1_n_547), .B
       (n_5988), .Q (n_6386));
  AND4X1 inc_add_1345_58_1_g866(.A (inc_add_1345_58_1_n_553), .B
       (n_5988), .C (n_6724), .D (n_4534), .Q
       (inc_add_1345_58_1_n_544));
  HAX1 inc_add_1345_58_1_g867(.A (inc_add_1345_58_1_n_550), .B
       (n_6724), .S (n_6388), .CO (inc_add_1345_58_1_n_547));
  HAX1 inc_add_1345_58_1_g868(.A (inc_add_1345_58_1_n_553), .B
       (n_4534), .S (n_6390), .CO (inc_add_1345_58_1_n_550));
  HAX1 inc_add_1345_58_1_g869(.A (inc_add_1345_58_1_n_556), .B
       (csr_mcycle[31]), .S (n_6392), .CO (inc_add_1345_58_1_n_553));
  EO2X1 inc_add_1345_58_1_g870(.A (inc_add_1345_58_1_n_559), .B
       (csr_mcycle[30]), .Q (n_6394));
  AND4X1 inc_add_1345_58_1_g871(.A (inc_add_1345_58_1_n_565), .B
       (csr_mcycle[28]), .C (csr_mcycle[29]), .D (csr_mcycle[30]), .Q
       (inc_add_1345_58_1_n_556));
  HAX1 inc_add_1345_58_1_g872(.A (inc_add_1345_58_1_n_562), .B
       (csr_mcycle[29]), .S (n_6396), .CO (inc_add_1345_58_1_n_559));
  HAX1 inc_add_1345_58_1_g873(.A (inc_add_1345_58_1_n_565), .B
       (csr_mcycle[28]), .S (n_6398), .CO (inc_add_1345_58_1_n_562));
  HAX1 inc_add_1345_58_1_g874(.A (inc_add_1345_58_1_n_568), .B
       (csr_mcycle[27]), .S (n_6400), .CO (inc_add_1345_58_1_n_565));
  EO2X1 inc_add_1345_58_1_g875(.A (inc_add_1345_58_1_n_573), .B
       (csr_mcycle[26]), .Q (n_6402));
  AND2X2 inc_add_1345_58_1_g876(.A (inc_add_1345_58_1_n_573), .B
       (csr_mcycle[26]), .Q (inc_add_1345_58_1_n_568));
  EO2X1 inc_add_1345_58_1_g877(.A (inc_add_1345_58_1_n_576), .B
       (csr_mcycle[25]), .Q (n_6404));
  AND4X1 inc_add_1345_58_1_g878(.A (inc_add_1345_58_1_n_582), .B
       (csr_mcycle[23]), .C (csr_mcycle[24]), .D (csr_mcycle[25]), .Q
       (inc_add_1345_58_1_n_573));
  HAX1 inc_add_1345_58_1_g879(.A (inc_add_1345_58_1_n_579), .B
       (csr_mcycle[24]), .S (n_6406), .CO (inc_add_1345_58_1_n_576));
  HAX1 inc_add_1345_58_1_g880(.A (inc_add_1345_58_1_n_582), .B
       (csr_mcycle[23]), .S (n_6408), .CO (inc_add_1345_58_1_n_579));
  HAX1 inc_add_1345_58_1_g881(.A (inc_add_1345_58_1_n_585), .B
       (csr_mcycle[22]), .S (n_6410), .CO (inc_add_1345_58_1_n_582));
  EO2X0 inc_add_1345_58_1_g882(.A (inc_add_1345_58_1_n_590), .B
       (csr_mcycle[21]), .Q (n_6412));
  AND2X2 inc_add_1345_58_1_g883(.A (inc_add_1345_58_1_n_590), .B
       (csr_mcycle[21]), .Q (inc_add_1345_58_1_n_585));
  EO2X0 inc_add_1345_58_1_g884(.A (inc_add_1345_58_1_n_595), .B
       (csr_mcycle[20]), .Q (n_6414));
  AND2X2 inc_add_1345_58_1_g885(.A (inc_add_1345_58_1_n_595), .B
       (csr_mcycle[20]), .Q (inc_add_1345_58_1_n_590));
  NO2I1X1 inc_add_1345_58_1_g887(.B (inc_add_1345_58_1_n_600), .AN
       (csr_mcycle[19]), .Q (inc_add_1345_58_1_n_595));
  EO2X0 inc_add_1345_58_1_g889(.A (inc_add_1345_58_1_n_605), .B
       (csr_mcycle[18]), .Q (n_6418));
  NA2X1 inc_add_1345_58_1_g890(.A (inc_add_1345_58_1_n_605), .B
       (csr_mcycle[18]), .Q (inc_add_1345_58_1_n_600));
  EO2X1 inc_add_1345_58_1_g891(.A (inc_add_1345_58_1_n_608), .B
       (csr_mcycle[17]), .Q (n_6420));
  AND4X1 inc_add_1345_58_1_g892(.A (inc_add_1345_58_1_n_614), .B
       (csr_mcycle[15]), .C (csr_mcycle[16]), .D (csr_mcycle[17]), .Q
       (inc_add_1345_58_1_n_605));
  HAX1 inc_add_1345_58_1_g893(.A (inc_add_1345_58_1_n_611), .B
       (csr_mcycle[16]), .S (n_6422), .CO (inc_add_1345_58_1_n_608));
  HAX1 inc_add_1345_58_1_g894(.A (inc_add_1345_58_1_n_614), .B
       (csr_mcycle[15]), .S (n_6424), .CO (inc_add_1345_58_1_n_611));
  HAX2 inc_add_1345_58_1_g895(.A (inc_add_1345_58_1_n_617), .B
       (csr_mcycle[14]), .S (n_6426), .CO (inc_add_1345_58_1_n_614));
  EO2X0 inc_add_1345_58_1_g896(.A (inc_add_1345_58_1_n_732), .B
       (csr_mcycle[13]), .Q (n_6428));
  AND2X2 inc_add_1345_58_1_g897(.A (inc_add_1345_58_1_n_732), .B
       (csr_mcycle[13]), .Q (inc_add_1345_58_1_n_617));
  EO2X0 inc_add_1345_58_1_g898(.A (inc_add_1345_58_1_n_627), .B
       (csr_mcycle[12]), .Q (n_6430));
  EO2X1 inc_add_1345_58_1_g901(.A (inc_add_1345_58_1_n_630), .B
       (csr_mcycle[11]), .Q (n_6432));
  AND4X1 inc_add_1345_58_1_g902(.A (inc_add_1345_58_1_n_638), .B
       (csr_mcycle[9]), .C (csr_mcycle[10]), .D (csr_mcycle[11]), .Q
       (inc_add_1345_58_1_n_627));
  HAX1 inc_add_1345_58_1_g903(.A (inc_add_1345_58_1_n_633), .B
       (csr_mcycle[10]), .S (n_6434), .CO (inc_add_1345_58_1_n_630));
  HAX1 inc_add_1345_58_1_g904(.A (inc_add_1345_58_1_n_638), .B
       (csr_mcycle[9]), .S (n_6436), .CO (inc_add_1345_58_1_n_633));
  EO2X1 inc_add_1345_58_1_g905(.A (inc_add_1345_58_1_n_643), .B
       (csr_mcycle[8]), .Q (n_6438));
  AND2X2 inc_add_1345_58_1_g906(.A (inc_add_1345_58_1_n_643), .B
       (csr_mcycle[8]), .Q (inc_add_1345_58_1_n_638));
  EO2X0 inc_add_1345_58_1_g907(.A (inc_add_1345_58_1_n_648), .B
       (csr_mcycle[7]), .Q (n_6440));
  AND2X4 inc_add_1345_58_1_g908(.A (inc_add_1345_58_1_n_648), .B
       (csr_mcycle[7]), .Q (inc_add_1345_58_1_n_643));
  NO2I1X1 inc_add_1345_58_1_g910(.B (inc_add_1345_58_1_n_653), .AN
       (csr_mcycle[6]), .Q (inc_add_1345_58_1_n_648));
  EO2X0 inc_add_1345_58_1_g912(.A (inc_add_1345_58_1_n_658), .B
       (csr_mcycle[5]), .Q (n_6444));
  NA2X1 inc_add_1345_58_1_g913(.A (inc_add_1345_58_1_n_658), .B
       (csr_mcycle[5]), .Q (inc_add_1345_58_1_n_653));
  NO2I1X1 inc_add_1345_58_1_g915(.B (inc_add_1345_58_1_n_663), .AN
       (csr_mcycle[4]), .Q (inc_add_1345_58_1_n_658));
  EO2X0 inc_add_1345_58_1_g917(.A (inc_add_1345_58_1_n_668), .B
       (csr_mcycle[3]), .Q (n_6448));
  NA2X1 inc_add_1345_58_1_g918(.A (inc_add_1345_58_1_n_668), .B
       (csr_mcycle[3]), .Q (inc_add_1345_58_1_n_663));
  NO2I1X1 inc_add_1345_58_1_g920(.B (inc_add_1345_58_1_n_673), .AN
       (csr_mcycle[2]), .Q (inc_add_1345_58_1_n_668));
  EO2X0 inc_add_1345_58_1_g922(.A (csr_mcycle[0]), .B (csr_mcycle[1]),
       .Q (n_6452));
  NA2X1 inc_add_1345_58_1_g923(.A (csr_mcycle[0]), .B (csr_mcycle[1]),
       .Q (inc_add_1345_58_1_n_673));
  EN2X0 inc_add_1345_58_1_g2(.A (inc_add_1345_58_1_n_471), .B (n_5737),
       .Q (n_6323));
  EN2X0 inc_add_1345_58_1_g926(.A (inc_add_1345_58_1_n_481), .B
       (n_5739), .Q (n_6346));
  AND2X1 inc_add_1345_58_1_g927(.A (inc_add_1345_58_1_n_494), .B
       (n_5742), .Q (inc_add_1345_58_1_n_728));
  EN2X0 inc_add_1345_58_1_g928(.A (inc_add_1345_58_1_n_504), .B
       (n_4536), .Q (n_6360));
  EN2X0 inc_add_1345_58_1_g929(.A (inc_add_1345_58_1_n_514), .B
       (n_5747), .Q (n_6364));
  EN2X1 inc_add_1345_58_1_g930(.A (inc_add_1345_58_1_n_600), .B
       (csr_mcycle[19]), .Q (n_6416));
  AND2X1 inc_add_1345_58_1_g931(.A (inc_add_1345_58_1_n_627), .B
       (csr_mcycle[12]), .Q (inc_add_1345_58_1_n_732));
  EN2X0 inc_add_1345_58_1_g932(.A (inc_add_1345_58_1_n_653), .B
       (csr_mcycle[6]), .Q (n_6442));
  EN2X0 inc_add_1345_58_1_g933(.A (inc_add_1345_58_1_n_663), .B
       (csr_mcycle[4]), .Q (n_6446));
  EN2X0 inc_add_1345_58_1_g934(.A (inc_add_1345_58_1_n_673), .B
       (csr_mcycle[2]), .Q (n_6450));
  EN2X1 inc_add_1345_58_1_g935(.A (inc_add_1345_58_1_n_448), .B
       (n_5985), .Q (n_6304));
  EO2X1 inc_add_1345_58_1_g936(.A (inc_add_1345_58_1_n_451), .B
       (n_5729), .Q (n_6306));
  NO2I1X2 inc_add_1345_58_1_g938(.B (inc_add_1345_58_1_n_514), .AN
       (n_5747), .Q (inc_add_1345_58_1_n_509));
  NA2X2 inc_add_1343_59_4_g1099(.A (inc_add_1343_59_4_n_708), .B
       (csr_mcycle[62]), .Q (inc_add_1343_59_4_n_703));
  MU2IX1 inc_add_1343_59_4_g1101(.S (inc_add_1343_59_4_n_713), .IN0
       (csr_mcycle[61]), .IN1 (inc_add_1343_59_4_n_1007), .Q (n_6242));
  NO2X4 inc_add_1343_59_4_g1102(.A (inc_add_1343_59_4_n_713), .B
       (inc_add_1343_59_4_n_1007), .Q (inc_add_1343_59_4_n_708));
  NA2X2 inc_add_1343_59_4_g1104(.A (inc_add_1343_59_4_n_718), .B
       (csr_mcycle[60]), .Q (inc_add_1343_59_4_n_713));
  MU2IX1 inc_add_1343_59_4_g1106(.S (inc_add_1343_59_4_n_724), .IN0
       (csr_mcycle[59]), .IN1 (inc_add_1343_59_4_n_972), .Q (n_6244));
  NO2X2 inc_add_1343_59_4_g1108(.A (inc_add_1343_59_4_n_724), .B
       (inc_add_1343_59_4_n_972), .Q (inc_add_1343_59_4_n_718));
  NA2X2 inc_add_1343_59_4_g1110(.A (inc_add_1343_59_4_n_727), .B
       (csr_mcycle[58]), .Q (inc_add_1343_59_4_n_724));
  MU2IX1 inc_add_1343_59_4_g1112(.S (inc_add_1343_59_4_n_735), .IN0
       (csr_mcycle[57]), .IN1 (inc_add_1343_59_4_n_968), .Q (n_6246));
  NO2X2 inc_add_1343_59_4_g1113(.A (inc_add_1343_59_4_n_735), .B
       (inc_add_1343_59_4_n_968), .Q (inc_add_1343_59_4_n_727));
  NA2X2 inc_add_1343_59_4_g1115(.A (inc_add_1343_59_4_n_740), .B
       (csr_mcycle[56]), .Q (inc_add_1343_59_4_n_735));
  AND6X2 inc_add_1343_59_4_g1119(.A (inc_add_1343_59_4_n_763), .B
       (csr_mcycle[51]), .C (csr_mcycle[53]), .D (csr_mcycle[52]), .E
       (csr_mcycle[54]), .F (csr_mcycle[55]), .Q
       (inc_add_1343_59_4_n_740));
  MU2IX1 inc_add_1343_59_4_g1120(.S (inc_add_1343_59_4_n_751), .IN0
       (csr_mcycle[54]), .IN1 (inc_add_1343_59_4_n_1010), .Q (n_6249));
  NO2X1 inc_add_1343_59_4_g1121(.A (inc_add_1343_59_4_n_751), .B
       (inc_add_1343_59_4_n_1010), .Q (inc_add_1343_59_4_n_745));
  NA2X1 inc_add_1343_59_4_g1123(.A (inc_add_1343_59_4_n_753), .B
       (csr_mcycle[53]), .Q (inc_add_1343_59_4_n_751));
  HAX2 inc_add_1343_59_4_g1125(.A (inc_add_1343_59_4_n_758), .B
       (csr_mcycle[52]), .S (n_6251), .CO (inc_add_1343_59_4_n_753));
  MU2IX1 inc_add_1343_59_4_g1126(.S (inc_add_1343_59_4_n_761), .IN0
       (csr_mcycle[51]), .IN1 (inc_add_1343_59_4_n_992), .Q (n_6252));
  NO2X1 inc_add_1343_59_4_g1127(.A (inc_add_1343_59_4_n_761), .B
       (inc_add_1343_59_4_n_992), .Q (inc_add_1343_59_4_n_758));
  INX1 inc_add_1343_59_4_g1129(.A (inc_add_1343_59_4_n_763), .Q
       (inc_add_1343_59_4_n_761));
  AND6X2 inc_add_1343_59_4_g1133(.A (inc_add_1343_59_4_n_783), .B
       (csr_mcycle[46]), .C (csr_mcycle[48]), .D (csr_mcycle[47]), .E
       (csr_mcycle[49]), .F (csr_mcycle[50]), .Q
       (inc_add_1343_59_4_n_763));
  NA2X1 inc_add_1343_59_4_g1135(.A (inc_add_1343_59_4_n_773), .B
       (csr_mcycle[49]), .Q (inc_add_1343_59_4_n_771));
  HAX2 inc_add_1343_59_4_g1137(.A (inc_add_1343_59_4_n_777), .B
       (csr_mcycle[48]), .S (n_6255), .CO (inc_add_1343_59_4_n_773));
  HAX2 inc_add_1343_59_4_g1138(.A (inc_add_1343_59_4_n_780), .B
       (csr_mcycle[47]), .S (n_6256), .CO (inc_add_1343_59_4_n_777));
  HAX2 inc_add_1343_59_4_g1139(.A (inc_add_1343_59_4_n_783), .B
       (csr_mcycle[46]), .S (n_6257), .CO (inc_add_1343_59_4_n_780));
  AND6X2 inc_add_1343_59_4_g1143(.A (inc_add_1343_59_4_n_805), .B
       (csr_mcycle[41]), .C (csr_mcycle[43]), .D (csr_mcycle[42]), .E
       (csr_mcycle[44]), .F (csr_mcycle[45]), .Q
       (inc_add_1343_59_4_n_783));
  NA2X1 inc_add_1343_59_4_g1145(.A (inc_add_1343_59_4_n_793), .B
       (csr_mcycle[44]), .Q (inc_add_1343_59_4_n_791));
  HAX2 inc_add_1343_59_4_g1147(.A (inc_add_1343_59_4_n_797), .B
       (csr_mcycle[43]), .S (n_6260), .CO (inc_add_1343_59_4_n_793));
  HAX2 inc_add_1343_59_4_g1148(.A (inc_add_1343_59_4_n_800), .B
       (csr_mcycle[42]), .S (n_6261), .CO (inc_add_1343_59_4_n_797));
  HAX2 inc_add_1343_59_4_g1149(.A (inc_add_1343_59_4_n_805), .B
       (csr_mcycle[41]), .S (n_6262), .CO (inc_add_1343_59_4_n_800));
  AND6X2 inc_add_1343_59_4_g1151(.A (inc_add_1343_59_4_n_824), .B
       (csr_mcycle[36]), .C (csr_mcycle[38]), .D (csr_mcycle[37]), .E
       (csr_mcycle[39]), .F (csr_mcycle[40]), .Q
       (inc_add_1343_59_4_n_805));
  NA2X1 inc_add_1343_59_4_g1153(.A (inc_add_1343_59_4_n_811), .B
       (csr_mcycle[39]), .Q (inc_add_1343_59_4_n_809));
  HAX2 inc_add_1343_59_4_g1155(.A (inc_add_1343_59_4_n_815), .B
       (csr_mcycle[38]), .S (n_6265), .CO (inc_add_1343_59_4_n_811));
  HAX2 inc_add_1343_59_4_g1156(.A (inc_add_1343_59_4_n_819), .B
       (csr_mcycle[37]), .S (n_6266), .CO (inc_add_1343_59_4_n_815));
  AND5X1 inc_add_1343_59_4_g1161(.A (inc_add_1343_59_4_n_835), .B
       (csr_mcycle[32]), .C (csr_mcycle[33]), .D (csr_mcycle[34]), .E
       (csr_mcycle[35]), .Q (inc_add_1343_59_4_n_824));
  HAX1 inc_add_1343_59_4_g1162(.A (inc_add_1343_59_4_n_832), .B
       (csr_mcycle[34]), .S (n_6269), .CO (inc_add_1343_59_4_n_830));
  HAX1 inc_add_1343_59_4_g1163(.A (inc_add_1343_59_4_n_834), .B
       (csr_mcycle[33]), .S (n_6270), .CO (inc_add_1343_59_4_n_832));
  HAX1 inc_add_1343_59_4_g1164(.A (inc_add_1343_59_4_n_835), .B
       (csr_mcycle[32]), .S (n_6271), .CO (inc_add_1343_59_4_n_834));
  EO2X1 inc_add_1343_59_4_g1166(.A (inc_add_1343_59_4_n_841), .B
       (n_5985), .Q (n_6272));
  AND6X2 inc_add_1343_59_4_g1167(.A (inc_add_1343_59_4_n_855), .B
       (n_5731), .C (n_5730), .D (n_5732), .E (n_5729), .F (n_5985), .Q
       (inc_add_1343_59_4_n_835));
  HAX1 inc_add_1343_59_4_g1168(.A (inc_add_1343_59_4_n_844), .B
       (n_5729), .S (n_6273), .CO (inc_add_1343_59_4_n_841));
  HAX1 inc_add_1343_59_4_g1169(.A (inc_add_1343_59_4_n_847), .B
       (n_5730), .S (n_6274), .CO (inc_add_1343_59_4_n_844));
  HAX1 inc_add_1343_59_4_g1170(.A (inc_add_1343_59_4_n_850), .B
       (n_5731), .S (n_6275), .CO (inc_add_1343_59_4_n_847));
  HAX1 inc_add_1343_59_4_g1171(.A (inc_add_1343_59_4_n_855), .B
       (n_5732), .S (n_6276), .CO (inc_add_1343_59_4_n_850));
  EO2X1 inc_add_1343_59_4_g1172(.A (inc_add_1343_59_4_n_858), .B
       (n_5733), .Q (n_6277));
  AND6X2 inc_add_1343_59_4_g1173(.A (inc_add_1343_59_4_n_870), .B
       (n_5737), .C (n_5736), .D (n_5735), .E (n_5734), .F (n_5733), .Q
       (inc_add_1343_59_4_n_855));
  HAX1 inc_add_1343_59_4_g1174(.A (inc_add_1343_59_4_n_861), .B
       (n_5734), .S (n_6278), .CO (inc_add_1343_59_4_n_858));
  HAX1 inc_add_1343_59_4_g1175(.A (inc_add_1343_59_4_n_864), .B
       (n_5735), .S (n_6279), .CO (inc_add_1343_59_4_n_861));
  HAX1 inc_add_1343_59_4_g1176(.A (inc_add_1343_59_4_n_867), .B
       (n_5736), .S (n_6280), .CO (inc_add_1343_59_4_n_864));
  HAX1 inc_add_1343_59_4_g1177(.A (inc_add_1343_59_4_n_870), .B
       (n_5737), .S (n_6281), .CO (inc_add_1343_59_4_n_867));
  HAX2 inc_add_1343_59_4_g1178(.A (inc_add_1343_59_4_n_873), .B
       (n_5738), .S (n_6282), .CO (inc_add_1343_59_4_n_870));
  EO2X1 inc_add_1343_59_4_g1179(.A (inc_add_1343_59_4_n_876), .B
       (n_5739), .Q (n_6283));
  AND5X2 inc_add_1343_59_4_g1180(.A (inc_add_1343_59_4_n_885), .B
       (n_5740), .C (n_5741), .D (n_5739), .E (n_5742), .Q
       (inc_add_1343_59_4_n_873));
  HAX1 inc_add_1343_59_4_g1181(.A (inc_add_1343_59_4_n_879), .B
       (n_5740), .S (n_6284), .CO (inc_add_1343_59_4_n_876));
  HAX1 inc_add_1343_59_4_g1182(.A (inc_add_1343_59_4_n_882), .B
       (n_5741), .S (n_6285), .CO (inc_add_1343_59_4_n_879));
  HAX1 inc_add_1343_59_4_g1183(.A (inc_add_1343_59_4_n_885), .B
       (n_5742), .S (n_6286), .CO (inc_add_1343_59_4_n_882));
  HAX1 inc_add_1343_59_4_g1184(.A (inc_add_1343_59_4_n_888), .B
       (n_5743), .S (n_6287), .CO (inc_add_1343_59_4_n_885));
  HAX1 inc_add_1343_59_4_g1185(.A (inc_add_1343_59_4_n_890), .B
       (n_4538), .S (n_6288), .CO (inc_add_1343_59_4_n_888));
  HAX1 inc_add_1343_59_4_g1186(.A (inc_add_1343_59_4_n_892), .B
       (n_4536), .S (n_6289), .CO (inc_add_1343_59_4_n_890));
  HAX1 inc_add_1343_59_4_g1187(.A (inc_add_1343_59_4_n_894), .B
       (n_5746), .S (n_6290), .CO (inc_add_1343_59_4_n_892));
  HAX2 inc_add_1343_59_4_g1188(.A (inc_add_1343_59_4_n_896), .B
       (n_5747), .S (n_6291), .CO (inc_add_1343_59_4_n_894));
  HAX2 inc_add_1343_59_4_g1189(.A (inc_add_1343_59_4_n_898), .B
       (n_5748), .S (n_6292), .CO (inc_add_1343_59_4_n_896));
  HAX2 inc_add_1343_59_4_g1190(.A (inc_add_1343_59_4_n_900), .B
       (n_5749), .S (n_6293), .CO (inc_add_1343_59_4_n_898));
  NO2I1X4 inc_add_1343_59_4_g1192(.B (inc_add_1343_59_4_n_905), .AN
       (n_5750), .Q (inc_add_1343_59_4_n_900));
  EO2X1 inc_add_1343_59_4_g1194(.A (inc_add_1343_59_4_n_911), .B
       (n_5751), .Q (n_6295));
  NA2X2 inc_add_1343_59_4_g1195(.A (inc_add_1343_59_4_n_911), .B
       (n_5751), .Q (inc_add_1343_59_4_n_905));
  EO2X1 inc_add_1343_59_4_g1197(.A (inc_add_1343_59_4_n_914), .B
       (n_4535), .Q (n_6299));
  NO2I1X1 inc_add_1343_59_4_g1198(.B (inc_add_1343_59_4_n_918), .AN
       (n_6726), .Q (inc_add_1343_59_4_n_911));
  HAX1 inc_add_1343_59_4_g1199(.A (inc_add_1343_59_4_n_923), .B
       (n_5987), .S (n_6300), .CO (inc_add_1343_59_4_n_914));
  EO2X1 inc_add_1343_59_4_g1201(.A (inc_add_1343_59_4_n_925), .B
       (n_6730), .Q (n_6297));
  NA2X2 inc_add_1343_59_4_g1202(.A (inc_add_1343_59_4_n_925), .B
       (n_6730), .Q (inc_add_1343_59_4_n_918));
  HAX1 inc_add_1343_59_4_g1203(.A (inc_add_1343_59_4_n_929), .B
       (n_5988), .S (n_6301), .CO (inc_add_1343_59_4_n_923));
  EO2X1 inc_add_1343_59_4_g1204(.A (inc_add_1343_59_4_n_930), .B
       (n_6731), .Q (n_6298));
  AND2X4 inc_add_1343_59_4_g1205(.A (inc_add_1343_59_4_n_930), .B
       (n_6731), .Q (inc_add_1343_59_4_n_925));
  HAX1 inc_add_1343_59_4_g1206(.A (n_6724), .B (n_4534), .S (n_6302),
       .CO (inc_add_1343_59_4_n_929));
  AND5X1 inc_add_1343_59_4_g1207(.A (n_5988), .B (n_4535), .C (n_6724),
       .D (n_4534), .E (n_5987), .Q (inc_add_1343_59_4_n_930));
  INX1 inc_add_1343_59_4_g1211(.A (csr_mcycle[57]), .Q
       (inc_add_1343_59_4_n_968));
  INX1 inc_add_1343_59_4_g1213(.A (csr_mcycle[59]), .Q
       (inc_add_1343_59_4_n_972));
  INX1 inc_add_1343_59_4_g1221(.A (csr_mcycle[51]), .Q
       (inc_add_1343_59_4_n_992));
  INX1 inc_add_1343_59_4_g1226(.A (csr_mcycle[61]), .Q
       (inc_add_1343_59_4_n_1007));
  INX1 inc_add_1343_59_4_g1227(.A (csr_mcycle[54]), .Q
       (inc_add_1343_59_4_n_1010));
  EO2X1 inc_add_1343_59_4_g2(.A (inc_add_1343_59_4_n_708), .B
       (csr_mcycle[62]), .Q (n_6241));
  EO2X1 inc_add_1343_59_4_g1228(.A (inc_add_1343_59_4_n_718), .B
       (csr_mcycle[60]), .Q (n_6243));
  EO2X1 inc_add_1343_59_4_g1229(.A (inc_add_1343_59_4_n_740), .B
       (csr_mcycle[56]), .Q (n_6247));
  EO2X1 inc_add_1343_59_4_g1230(.A (inc_add_1343_59_4_n_753), .B
       (csr_mcycle[53]), .Q (n_6250));
  EO2X1 inc_add_1343_59_4_g1231(.A (inc_add_1343_59_4_n_773), .B
       (csr_mcycle[49]), .Q (n_6254));
  EO2X1 inc_add_1343_59_4_g1232(.A (inc_add_1343_59_4_n_793), .B
       (csr_mcycle[44]), .Q (n_6259));
  EO2X1 inc_add_1343_59_4_g1233(.A (inc_add_1343_59_4_n_811), .B
       (csr_mcycle[39]), .Q (n_6264));
  EO2X1 inc_add_1343_59_4_g1234(.A (inc_add_1343_59_4_n_824), .B
       (csr_mcycle[36]), .Q (n_6267));
  EN2X1 inc_add_1343_59_4_g1235(.A (inc_add_1343_59_4_n_905), .B
       (n_5750), .Q (n_6294));
  EN2X1 inc_add_1343_59_4_g1236(.A (inc_add_1343_59_4_n_918), .B
       (n_6726), .Q (n_6296));
  EN2X1 inc_add_1343_59_4_g1237(.A (inc_add_1343_59_4_n_703), .B
       (csr_mcycle[63]), .Q (n_6240));
  EO2X1 inc_add_1343_59_4_g1238(.A (inc_add_1343_59_4_n_745), .B
       (csr_mcycle[55]), .Q (n_6248));
  EN2X1 inc_add_1343_59_4_g1239(.A (inc_add_1343_59_4_n_771), .B
       (csr_mcycle[50]), .Q (n_6253));
  EN2X1 inc_add_1343_59_4_g1240(.A (inc_add_1343_59_4_n_809), .B
       (csr_mcycle[40]), .Q (n_6263));
  EN2X1 inc_add_1343_59_4_g1241(.A (inc_add_1343_59_4_n_791), .B
       (csr_mcycle[45]), .Q (n_6258));
  EO2X1 inc_add_1343_59_4_g1242(.A (inc_add_1343_59_4_n_727), .B
       (csr_mcycle[58]), .Q (n_6245));
  EO2X1 inc_add_1343_59_4_g1243(.A (inc_add_1343_59_4_n_830), .B
       (csr_mcycle[35]), .Q (n_6268));
  AND6X1 inc_add_1343_59_4_g1245(.A (inc_add_1343_59_4_n_835), .B
       (csr_mcycle[32]), .C (csr_mcycle[34]), .D (csr_mcycle[33]), .E
       (csr_mcycle[35]), .F (csr_mcycle[36]), .Q
       (inc_add_1343_59_4_n_819));
  NA2X1 inc_add_1347_34_2_g819(.A (inc_add_1347_34_2_n_451), .B
       (csr_mcycle[62]), .Q (inc_add_1347_34_2_n_448));
  HAX2 inc_add_1347_34_2_g820(.A (inc_add_1347_34_2_n_454), .B
       (csr_mcycle[61]), .S (n_6307), .CO (inc_add_1347_34_2_n_451));
  HAX2 inc_add_1347_34_2_g821(.A (inc_add_1347_34_2_n_456), .B
       (csr_mcycle[60]), .S (n_6309), .CO (inc_add_1347_34_2_n_454));
  HAX2 inc_add_1347_34_2_g822(.A (inc_add_1347_34_2_n_458), .B
       (csr_mcycle[59]), .S (n_6311), .CO (inc_add_1347_34_2_n_456));
  HAX2 inc_add_1347_34_2_g823(.A (inc_add_1347_34_2_n_460), .B
       (csr_mcycle[58]), .S (n_6313), .CO (inc_add_1347_34_2_n_458));
  HAX2 inc_add_1347_34_2_g824(.A (inc_add_1347_34_2_n_462), .B
       (csr_mcycle[57]), .S (n_6315), .CO (inc_add_1347_34_2_n_460));
  HAX2 inc_add_1347_34_2_g825(.A (inc_add_1347_34_2_n_464), .B
       (csr_mcycle[56]), .S (n_6317), .CO (inc_add_1347_34_2_n_462));
  HAX2 inc_add_1347_34_2_g826(.A (inc_add_1347_34_2_n_466), .B
       (csr_mcycle[55]), .S (n_6319), .CO (inc_add_1347_34_2_n_464));
  HAX2 inc_add_1347_34_2_g827(.A (inc_add_1347_34_2_n_468), .B
       (csr_mcycle[54]), .S (n_6321), .CO (inc_add_1347_34_2_n_466));
  HAX2 inc_add_1347_34_2_g828(.A (inc_add_1347_34_2_n_470), .B
       (csr_mcycle[53]), .S (n_6329), .CO (inc_add_1347_34_2_n_468));
  HAX2 inc_add_1347_34_2_g829(.A (inc_add_1347_34_2_n_472), .B
       (csr_mcycle[52]), .S (n_6341), .CO (inc_add_1347_34_2_n_470));
  HAX2 inc_add_1347_34_2_g830(.A (inc_add_1347_34_2_n_474), .B
       (csr_mcycle[51]), .S (n_6349), .CO (inc_add_1347_34_2_n_472));
  EO2X0 inc_add_1347_34_2_g834(.A (inc_add_1347_34_2_n_484), .B
       (csr_mcycle[49]), .Q (n_6353));
  NA2X1 inc_add_1347_34_2_g835(.A (inc_add_1347_34_2_n_484), .B
       (csr_mcycle[49]), .Q (inc_add_1347_34_2_n_479));
  NO2I1X4 inc_add_1347_34_2_g837(.B (inc_add_1347_34_2_n_489), .AN
       (csr_mcycle[48]), .Q (inc_add_1347_34_2_n_484));
  EO2X0 inc_add_1347_34_2_g839(.A (inc_add_1347_34_2_n_494), .B
       (csr_mcycle[47]), .Q (n_6357));
  NA2X4 inc_add_1347_34_2_g840(.A (inc_add_1347_34_2_n_494), .B
       (csr_mcycle[47]), .Q (inc_add_1347_34_2_n_489));
  EO2X0 inc_add_1347_34_2_g844(.A (inc_add_1347_34_2_n_504), .B
       (csr_mcycle[45]), .Q (n_6361));
  NA2X2 inc_add_1347_34_2_g845(.A (inc_add_1347_34_2_n_504), .B
       (csr_mcycle[45]), .Q (inc_add_1347_34_2_n_499));
  EO2X0 inc_add_1347_34_2_g846(.A (inc_add_1347_34_2_n_509), .B
       (csr_mcycle[44]), .Q (n_6363));
  AND2X4 inc_add_1347_34_2_g847(.A (inc_add_1347_34_2_n_509), .B
       (csr_mcycle[44]), .Q (inc_add_1347_34_2_n_504));
  EO2X0 inc_add_1347_34_2_g848(.A (inc_add_1347_34_2_n_514), .B
       (csr_mcycle[43]), .Q (n_6365));
  AND2X1 inc_add_1347_34_2_g849(.A (inc_add_1347_34_2_n_514), .B
       (csr_mcycle[43]), .Q (inc_add_1347_34_2_n_509));
  EO2X0 inc_add_1347_34_2_g850(.A (inc_add_1347_34_2_n_517), .B
       (csr_mcycle[42]), .Q (n_6368));
  AND2X1 inc_add_1347_34_2_g851(.A (inc_add_1347_34_2_n_517), .B
       (csr_mcycle[42]), .Q (inc_add_1347_34_2_n_514));
  HAX2 inc_add_1347_34_2_g852(.A (inc_add_1347_34_2_n_520), .B
       (csr_mcycle[41]), .S (n_6370), .CO (inc_add_1347_34_2_n_517));
  EO2X1 inc_add_1347_34_2_g853(.A (inc_add_1347_34_2_n_523), .B
       (csr_mcycle[40]), .Q (n_6372));
  AND3X1 inc_add_1347_34_2_g854(.A (inc_add_1347_34_2_n_526), .B
       (csr_mcycle[39]), .C (csr_mcycle[40]), .Q
       (inc_add_1347_34_2_n_520));
  HAX1 inc_add_1347_34_2_g855(.A (inc_add_1347_34_2_n_526), .B
       (csr_mcycle[39]), .S (n_6375), .CO (inc_add_1347_34_2_n_523));
  HAX2 inc_add_1347_34_2_g856(.A (inc_add_1347_34_2_n_529), .B
       (csr_mcycle[38]), .S (n_6377), .CO (inc_add_1347_34_2_n_526));
  EO2X1 inc_add_1347_34_2_g857(.A (inc_add_1347_34_2_n_532), .B
       (csr_mcycle[37]), .Q (n_6379));
  AND4X1 inc_add_1347_34_2_g858(.A (inc_add_1347_34_2_n_538), .B
       (csr_mcycle[35]), .C (csr_mcycle[36]), .D (csr_mcycle[37]), .Q
       (inc_add_1347_34_2_n_529));
  HAX1 inc_add_1347_34_2_g859(.A (inc_add_1347_34_2_n_535), .B
       (csr_mcycle[36]), .S (n_6381), .CO (inc_add_1347_34_2_n_532));
  HAX1 inc_add_1347_34_2_g860(.A (inc_add_1347_34_2_n_538), .B
       (csr_mcycle[35]), .S (n_6383), .CO (inc_add_1347_34_2_n_535));
  HAX1 inc_add_1347_34_2_g861(.A (inc_add_1347_34_2_n_541), .B
       (csr_mcycle[34]), .S (n_6385), .CO (inc_add_1347_34_2_n_538));
  EO2X0 inc_add_1347_34_2_g862(.A (inc_add_1347_34_2_n_546), .B
       (csr_mcycle[33]), .Q (n_6387));
  AND2X2 inc_add_1347_34_2_g863(.A (inc_add_1347_34_2_n_546), .B
       (csr_mcycle[33]), .Q (inc_add_1347_34_2_n_541));
  EO2X1 inc_add_1347_34_2_g864(.A (inc_add_1347_34_2_n_549), .B
       (csr_mcycle[32]), .Q (n_6389));
  AND4X1 inc_add_1347_34_2_g865(.A (inc_add_1347_34_2_n_555), .B
       (csr_mcycle[30]), .C (csr_mcycle[31]), .D (csr_mcycle[32]), .Q
       (inc_add_1347_34_2_n_546));
  HAX1 inc_add_1347_34_2_g866(.A (inc_add_1347_34_2_n_552), .B
       (csr_mcycle[31]), .S (n_6391), .CO (inc_add_1347_34_2_n_549));
  HAX1 inc_add_1347_34_2_g867(.A (inc_add_1347_34_2_n_555), .B
       (csr_mcycle[30]), .S (n_6393), .CO (inc_add_1347_34_2_n_552));
  HAX1 inc_add_1347_34_2_g868(.A (inc_add_1347_34_2_n_558), .B
       (csr_mcycle[29]), .S (n_6395), .CO (inc_add_1347_34_2_n_555));
  NO2I1X1 inc_add_1347_34_2_g870(.B (inc_add_1347_34_2_n_563), .AN
       (csr_mcycle[28]), .Q (inc_add_1347_34_2_n_558));
  EO2X0 inc_add_1347_34_2_g872(.A (inc_add_1347_34_2_n_568), .B
       (csr_mcycle[27]), .Q (n_6399));
  NA2X1 inc_add_1347_34_2_g873(.A (inc_add_1347_34_2_n_568), .B
       (csr_mcycle[27]), .Q (inc_add_1347_34_2_n_563));
  EO2X1 inc_add_1347_34_2_g874(.A (inc_add_1347_34_2_n_571), .B
       (csr_mcycle[26]), .Q (n_6401));
  AND4X1 inc_add_1347_34_2_g875(.A (inc_add_1347_34_2_n_577), .B
       (csr_mcycle[24]), .C (csr_mcycle[25]), .D (csr_mcycle[26]), .Q
       (inc_add_1347_34_2_n_568));
  HAX1 inc_add_1347_34_2_g876(.A (inc_add_1347_34_2_n_574), .B
       (csr_mcycle[25]), .S (n_6403), .CO (inc_add_1347_34_2_n_571));
  HAX1 inc_add_1347_34_2_g877(.A (inc_add_1347_34_2_n_577), .B
       (csr_mcycle[24]), .S (n_6405), .CO (inc_add_1347_34_2_n_574));
  HAX2 inc_add_1347_34_2_g878(.A (inc_add_1347_34_2_n_580), .B
       (csr_mcycle[23]), .S (n_6407), .CO (inc_add_1347_34_2_n_577));
  EO2X0 inc_add_1347_34_2_g879(.A (inc_add_1347_34_2_n_585), .B
       (csr_mcycle[22]), .Q (n_6409));
  AND2X2 inc_add_1347_34_2_g880(.A (inc_add_1347_34_2_n_585), .B
       (csr_mcycle[22]), .Q (inc_add_1347_34_2_n_580));
  NO2I1X1 inc_add_1347_34_2_g882(.B (inc_add_1347_34_2_n_590), .AN
       (csr_mcycle[21]), .Q (inc_add_1347_34_2_n_585));
  EO2X0 inc_add_1347_34_2_g884(.A (inc_add_1347_34_2_n_595), .B
       (csr_mcycle[20]), .Q (n_6413));
  NA2X1 inc_add_1347_34_2_g885(.A (inc_add_1347_34_2_n_595), .B
       (csr_mcycle[20]), .Q (inc_add_1347_34_2_n_590));
  EO2X1 inc_add_1347_34_2_g886(.A (inc_add_1347_34_2_n_598), .B
       (csr_mcycle[19]), .Q (n_6415));
  AND4X1 inc_add_1347_34_2_g887(.A (inc_add_1347_34_2_n_604), .B
       (csr_mcycle[17]), .C (csr_mcycle[18]), .D (csr_mcycle[19]), .Q
       (inc_add_1347_34_2_n_595));
  HAX1 inc_add_1347_34_2_g888(.A (inc_add_1347_34_2_n_601), .B
       (csr_mcycle[18]), .S (n_6417), .CO (inc_add_1347_34_2_n_598));
  HAX1 inc_add_1347_34_2_g889(.A (inc_add_1347_34_2_n_604), .B
       (csr_mcycle[17]), .S (n_6419), .CO (inc_add_1347_34_2_n_601));
  HAX2 inc_add_1347_34_2_g890(.A (inc_add_1347_34_2_n_607), .B
       (csr_mcycle[16]), .S (n_6421), .CO (inc_add_1347_34_2_n_604));
  NO2I1X1 inc_add_1347_34_2_g892(.B (inc_add_1347_34_2_n_612), .AN
       (csr_mcycle[15]), .Q (inc_add_1347_34_2_n_607));
  EO2X0 inc_add_1347_34_2_g894(.A (inc_add_1347_34_2_n_617), .B
       (csr_mcycle[14]), .Q (n_6425));
  NA2X1 inc_add_1347_34_2_g895(.A (inc_add_1347_34_2_n_617), .B
       (csr_mcycle[14]), .Q (inc_add_1347_34_2_n_612));
  EO2X1 inc_add_1347_34_2_g896(.A (inc_add_1347_34_2_n_620), .B
       (csr_mcycle[13]), .Q (n_6427));
  AND4X1 inc_add_1347_34_2_g897(.A (inc_add_1347_34_2_n_626), .B
       (csr_mcycle[11]), .C (csr_mcycle[12]), .D (csr_mcycle[13]), .Q
       (inc_add_1347_34_2_n_617));
  HAX1 inc_add_1347_34_2_g898(.A (inc_add_1347_34_2_n_623), .B
       (csr_mcycle[12]), .S (n_6429), .CO (inc_add_1347_34_2_n_620));
  HAX1 inc_add_1347_34_2_g899(.A (inc_add_1347_34_2_n_626), .B
       (csr_mcycle[11]), .S (n_6431), .CO (inc_add_1347_34_2_n_623));
  HAX2 inc_add_1347_34_2_g900(.A (inc_add_1347_34_2_n_629), .B
       (csr_mcycle[10]), .S (n_6433), .CO (inc_add_1347_34_2_n_626));
  EO2X0 inc_add_1347_34_2_g901(.A (inc_add_1347_34_2_n_634), .B
       (csr_mcycle[9]), .Q (n_6435));
  AND2X2 inc_add_1347_34_2_g902(.A (inc_add_1347_34_2_n_634), .B
       (csr_mcycle[9]), .Q (inc_add_1347_34_2_n_629));
  NO2I1X1 inc_add_1347_34_2_g904(.B (inc_add_1347_34_2_n_639), .AN
       (csr_mcycle[8]), .Q (inc_add_1347_34_2_n_634));
  EO2X0 inc_add_1347_34_2_g906(.A (inc_add_1347_34_2_n_644), .B
       (csr_mcycle[7]), .Q (n_6439));
  NA2X2 inc_add_1347_34_2_g907(.A (inc_add_1347_34_2_n_644), .B
       (csr_mcycle[7]), .Q (inc_add_1347_34_2_n_639));
  NO2I1X2 inc_add_1347_34_2_g909(.B (inc_add_1347_34_2_n_649), .AN
       (csr_mcycle[6]), .Q (inc_add_1347_34_2_n_644));
  EO2X0 inc_add_1347_34_2_g911(.A (inc_add_1347_34_2_n_654), .B
       (csr_mcycle[5]), .Q (n_6443));
  NA2X2 inc_add_1347_34_2_g912(.A (inc_add_1347_34_2_n_654), .B
       (csr_mcycle[5]), .Q (inc_add_1347_34_2_n_649));
  NO2I1X1 inc_add_1347_34_2_g914(.B (inc_add_1347_34_2_n_659), .AN
       (csr_mcycle[4]), .Q (inc_add_1347_34_2_n_654));
  EO2X0 inc_add_1347_34_2_g916(.A (inc_add_1347_34_2_n_664), .B
       (csr_mcycle[3]), .Q (n_6447));
  NA2X2 inc_add_1347_34_2_g917(.A (inc_add_1347_34_2_n_664), .B
       (csr_mcycle[3]), .Q (inc_add_1347_34_2_n_659));
  NO2I1X1 inc_add_1347_34_2_g919(.B (inc_add_1347_34_2_n_669), .AN
       (csr_mcycle[2]), .Q (inc_add_1347_34_2_n_664));
  EO2X0 inc_add_1347_34_2_g921(.A (csr_mcycle[0]), .B (csr_mcycle[1]),
       .Q (n_6451));
  NA2X1 inc_add_1347_34_2_g922(.A (csr_mcycle[0]), .B (csr_mcycle[1]),
       .Q (inc_add_1347_34_2_n_669));
  EN2X0 inc_add_1347_34_2_g2(.A (inc_add_1347_34_2_n_479), .B
       (csr_mcycle[50]), .Q (n_6351));
  EN2X0 inc_add_1347_34_2_g925(.A (inc_add_1347_34_2_n_489), .B
       (csr_mcycle[48]), .Q (n_6355));
  EN2X0 inc_add_1347_34_2_g926(.A (inc_add_1347_34_2_n_499), .B
       (csr_mcycle[46]), .Q (n_6359));
  EN2X1 inc_add_1347_34_2_g927(.A (inc_add_1347_34_2_n_563), .B
       (csr_mcycle[28]), .Q (n_6397));
  EN2X1 inc_add_1347_34_2_g928(.A (inc_add_1347_34_2_n_590), .B
       (csr_mcycle[21]), .Q (n_6411));
  EN2X1 inc_add_1347_34_2_g929(.A (inc_add_1347_34_2_n_612), .B
       (csr_mcycle[15]), .Q (n_6423));
  EN2X0 inc_add_1347_34_2_g930(.A (inc_add_1347_34_2_n_639), .B
       (csr_mcycle[8]), .Q (n_6437));
  EN2X0 inc_add_1347_34_2_g931(.A (inc_add_1347_34_2_n_649), .B
       (csr_mcycle[6]), .Q (n_6441));
  EN2X0 inc_add_1347_34_2_g932(.A (inc_add_1347_34_2_n_659), .B
       (csr_mcycle[4]), .Q (n_6445));
  EN2X0 inc_add_1347_34_2_g933(.A (inc_add_1347_34_2_n_669), .B
       (csr_mcycle[2]), .Q (n_6449));
  EN2X1 inc_add_1347_34_2_g934(.A (inc_add_1347_34_2_n_448), .B
       (csr_mcycle[63]), .Q (n_6303));
  EO2X1 inc_add_1347_34_2_g935(.A (inc_add_1347_34_2_n_451), .B
       (csr_mcycle[62]), .Q (n_6305));
  NO2I1X1 inc_add_1347_34_2_g937(.B (inc_add_1347_34_2_n_479), .AN
       (csr_mcycle[50]), .Q (inc_add_1347_34_2_n_474));
  NO2I1X2 inc_add_1347_34_2_g939(.B (inc_add_1347_34_2_n_499), .AN
       (csr_mcycle[46]), .Q (inc_add_1347_34_2_n_494));
  NA2X2 inc_ADD_UNS_OP5494_3_g829(.A (inc_ADD_UNS_OP5494_3_n_455), .B
       (csr_minstret[62]), .Q (inc_ADD_UNS_OP5494_3_n_452));
  HAX2 inc_ADD_UNS_OP5494_3_g831(.A (inc_ADD_UNS_OP5494_3_n_458), .B
       (csr_minstret[61]), .S (n_5823), .CO
       (inc_ADD_UNS_OP5494_3_n_455));
  HAX2 inc_ADD_UNS_OP5494_3_g832(.A (inc_ADD_UNS_OP5494_3_n_460), .B
       (csr_minstret[60]), .S (n_5825), .CO
       (inc_ADD_UNS_OP5494_3_n_458));
  HAX2 inc_ADD_UNS_OP5494_3_g833(.A (inc_ADD_UNS_OP5494_3_n_462), .B
       (csr_minstret[59]), .S (n_5827), .CO
       (inc_ADD_UNS_OP5494_3_n_460));
  HAX2 inc_ADD_UNS_OP5494_3_g834(.A (inc_ADD_UNS_OP5494_3_n_464), .B
       (csr_minstret[58]), .S (n_5829), .CO
       (inc_ADD_UNS_OP5494_3_n_462));
  HAX2 inc_ADD_UNS_OP5494_3_g835(.A (inc_ADD_UNS_OP5494_3_n_466), .B
       (csr_minstret[57]), .S (n_5831), .CO
       (inc_ADD_UNS_OP5494_3_n_464));
  HAX2 inc_ADD_UNS_OP5494_3_g836(.A (inc_ADD_UNS_OP5494_3_n_468), .B
       (csr_minstret[56]), .S (n_5833), .CO
       (inc_ADD_UNS_OP5494_3_n_466));
  HAX2 inc_ADD_UNS_OP5494_3_g837(.A (inc_ADD_UNS_OP5494_3_n_470), .B
       (csr_minstret[55]), .S (n_5835), .CO
       (inc_ADD_UNS_OP5494_3_n_468));
  HAX2 inc_ADD_UNS_OP5494_3_g838(.A (inc_ADD_UNS_OP5494_3_n_472), .B
       (csr_minstret[54]), .S (n_5837), .CO
       (inc_ADD_UNS_OP5494_3_n_470));
  HAX2 inc_ADD_UNS_OP5494_3_g839(.A (inc_ADD_UNS_OP5494_3_n_474), .B
       (csr_minstret[53]), .S (n_5839), .CO
       (inc_ADD_UNS_OP5494_3_n_472));
  HAX2 inc_ADD_UNS_OP5494_3_g840(.A (inc_ADD_UNS_OP5494_3_n_476), .B
       (csr_minstret[52]), .S (n_5841), .CO
       (inc_ADD_UNS_OP5494_3_n_474));
  HAX2 inc_ADD_UNS_OP5494_3_g841(.A (inc_ADD_UNS_OP5494_3_n_478), .B
       (csr_minstret[51]), .S (n_5843), .CO
       (inc_ADD_UNS_OP5494_3_n_476));
  EO2X0 inc_ADD_UNS_OP5494_3_g845(.A (inc_ADD_UNS_OP5494_3_n_488), .B
       (csr_minstret[49]), .Q (n_5847));
  NA2X2 inc_ADD_UNS_OP5494_3_g846(.A (inc_ADD_UNS_OP5494_3_n_488), .B
       (csr_minstret[49]), .Q (inc_ADD_UNS_OP5494_3_n_483));
  NO2I1X4 inc_ADD_UNS_OP5494_3_g848(.B (inc_ADD_UNS_OP5494_3_n_493),
       .AN (csr_minstret[48]), .Q (inc_ADD_UNS_OP5494_3_n_488));
  EO2X0 inc_ADD_UNS_OP5494_3_g850(.A (inc_ADD_UNS_OP5494_3_n_498), .B
       (csr_minstret[47]), .Q (n_5851));
  NA2X2 inc_ADD_UNS_OP5494_3_g851(.A (inc_ADD_UNS_OP5494_3_n_498), .B
       (csr_minstret[47]), .Q (inc_ADD_UNS_OP5494_3_n_493));
  NO2I1X4 inc_ADD_UNS_OP5494_3_g853(.B (inc_ADD_UNS_OP5494_3_n_503),
       .AN (csr_minstret[46]), .Q (inc_ADD_UNS_OP5494_3_n_498));
  EO2X0 inc_ADD_UNS_OP5494_3_g855(.A (inc_ADD_UNS_OP5494_3_n_508), .B
       (csr_minstret[45]), .Q (n_5855));
  NA2X2 inc_ADD_UNS_OP5494_3_g856(.A (inc_ADD_UNS_OP5494_3_n_508), .B
       (csr_minstret[45]), .Q (inc_ADD_UNS_OP5494_3_n_503));
  NO2I1X4 inc_ADD_UNS_OP5494_3_g858(.B (inc_ADD_UNS_OP5494_3_n_513),
       .AN (csr_minstret[44]), .Q (inc_ADD_UNS_OP5494_3_n_508));
  EO2X0 inc_ADD_UNS_OP5494_3_g860(.A (inc_ADD_UNS_OP5494_3_n_518), .B
       (csr_minstret[43]), .Q (n_5859));
  NA2X2 inc_ADD_UNS_OP5494_3_g861(.A (inc_ADD_UNS_OP5494_3_n_518), .B
       (csr_minstret[43]), .Q (inc_ADD_UNS_OP5494_3_n_513));
  EO2X1 inc_ADD_UNS_OP5494_3_g862(.A (inc_ADD_UNS_OP5494_3_n_521), .B
       (csr_minstret[42]), .Q (n_5861));
  AND6X2 inc_ADD_UNS_OP5494_3_g863(.A (inc_ADD_UNS_OP5494_3_n_533), .B
       (csr_minstret[38]), .C (csr_minstret[40]), .D
       (csr_minstret[39]), .E (csr_minstret[41]), .F
       (csr_minstret[42]), .Q (inc_ADD_UNS_OP5494_3_n_518));
  HAX1 inc_ADD_UNS_OP5494_3_g864(.A (inc_ADD_UNS_OP5494_3_n_524), .B
       (csr_minstret[41]), .S (n_5863), .CO
       (inc_ADD_UNS_OP5494_3_n_521));
  HAX1 inc_ADD_UNS_OP5494_3_g865(.A (inc_ADD_UNS_OP5494_3_n_527), .B
       (csr_minstret[40]), .S (n_5865), .CO
       (inc_ADD_UNS_OP5494_3_n_524));
  HAX1 inc_ADD_UNS_OP5494_3_g866(.A (inc_ADD_UNS_OP5494_3_n_530), .B
       (csr_minstret[39]), .S (n_5867), .CO
       (inc_ADD_UNS_OP5494_3_n_527));
  HAX1 inc_ADD_UNS_OP5494_3_g867(.A (inc_ADD_UNS_OP5494_3_n_533), .B
       (csr_minstret[38]), .S (n_5869), .CO
       (inc_ADD_UNS_OP5494_3_n_530));
  HAX2 inc_ADD_UNS_OP5494_3_g868(.A (inc_ADD_UNS_OP5494_3_n_536), .B
       (csr_minstret[37]), .S (n_5871), .CO
       (inc_ADD_UNS_OP5494_3_n_533));
  EO2X1 inc_ADD_UNS_OP5494_3_g869(.A (inc_ADD_UNS_OP5494_3_n_539), .B
       (csr_minstret[36]), .Q (n_5873));
  AND3X1 inc_ADD_UNS_OP5494_3_g870(.A (inc_ADD_UNS_OP5494_3_n_542), .B
       (csr_minstret[35]), .C (csr_minstret[36]), .Q
       (inc_ADD_UNS_OP5494_3_n_536));
  HAX1 inc_ADD_UNS_OP5494_3_g871(.A (inc_ADD_UNS_OP5494_3_n_542), .B
       (csr_minstret[35]), .S (n_5875), .CO
       (inc_ADD_UNS_OP5494_3_n_539));
  HAX2 inc_ADD_UNS_OP5494_3_g872(.A (inc_ADD_UNS_OP5494_3_n_545), .B
       (csr_minstret[34]), .S (n_5877), .CO
       (inc_ADD_UNS_OP5494_3_n_542));
  EO2X1 inc_ADD_UNS_OP5494_3_g873(.A (inc_ADD_UNS_OP5494_3_n_548), .B
       (csr_minstret[33]), .Q (n_5879));
  AND4X1 inc_ADD_UNS_OP5494_3_g874(.A (inc_ADD_UNS_OP5494_3_n_554), .B
       (csr_minstret[31]), .C (csr_minstret[32]), .D
       (csr_minstret[33]), .Q (inc_ADD_UNS_OP5494_3_n_545));
  HAX1 inc_ADD_UNS_OP5494_3_g875(.A (inc_ADD_UNS_OP5494_3_n_551), .B
       (csr_minstret[32]), .S (n_5881), .CO
       (inc_ADD_UNS_OP5494_3_n_548));
  HAX1 inc_ADD_UNS_OP5494_3_g876(.A (inc_ADD_UNS_OP5494_3_n_554), .B
       (csr_minstret[31]), .S (n_5883), .CO
       (inc_ADD_UNS_OP5494_3_n_551));
  HAX1 inc_ADD_UNS_OP5494_3_g877(.A (inc_ADD_UNS_OP5494_3_n_557), .B
       (csr_minstret[30]), .S (n_5885), .CO
       (inc_ADD_UNS_OP5494_3_n_554));
  EO2X0 inc_ADD_UNS_OP5494_3_g878(.A (inc_ADD_UNS_OP5494_3_n_562), .B
       (csr_minstret[29]), .Q (n_5887));
  AND2X2 inc_ADD_UNS_OP5494_3_g879(.A (inc_ADD_UNS_OP5494_3_n_562), .B
       (csr_minstret[29]), .Q (inc_ADD_UNS_OP5494_3_n_557));
  EO2X0 inc_ADD_UNS_OP5494_3_g880(.A (inc_ADD_UNS_OP5494_3_n_567), .B
       (csr_minstret[28]), .Q (n_5889));
  AND2X2 inc_ADD_UNS_OP5494_3_g881(.A (inc_ADD_UNS_OP5494_3_n_567), .B
       (csr_minstret[28]), .Q (inc_ADD_UNS_OP5494_3_n_562));
  NO2I1X1 inc_ADD_UNS_OP5494_3_g883(.B (inc_ADD_UNS_OP5494_3_n_572),
       .AN (csr_minstret[27]), .Q (inc_ADD_UNS_OP5494_3_n_567));
  EO2X0 inc_ADD_UNS_OP5494_3_g885(.A (inc_ADD_UNS_OP5494_3_n_577), .B
       (csr_minstret[26]), .Q (n_5893));
  NA2X1 inc_ADD_UNS_OP5494_3_g886(.A (inc_ADD_UNS_OP5494_3_n_577), .B
       (csr_minstret[26]), .Q (inc_ADD_UNS_OP5494_3_n_572));
  EO2X0 inc_ADD_UNS_OP5494_3_g887(.A (inc_ADD_UNS_OP5494_3_n_582), .B
       (csr_minstret[25]), .Q (n_5895));
  AND2X2 inc_ADD_UNS_OP5494_3_g888(.A (inc_ADD_UNS_OP5494_3_n_582), .B
       (csr_minstret[25]), .Q (inc_ADD_UNS_OP5494_3_n_577));
  EO2X1 inc_ADD_UNS_OP5494_3_g889(.A (inc_ADD_UNS_OP5494_3_n_585), .B
       (csr_minstret[24]), .Q (n_5897));
  AND4X1 inc_ADD_UNS_OP5494_3_g890(.A (inc_ADD_UNS_OP5494_3_n_591), .B
       (csr_minstret[22]), .C (csr_minstret[23]), .D
       (csr_minstret[24]), .Q (inc_ADD_UNS_OP5494_3_n_582));
  HAX1 inc_ADD_UNS_OP5494_3_g891(.A (inc_ADD_UNS_OP5494_3_n_588), .B
       (csr_minstret[23]), .S (n_5899), .CO
       (inc_ADD_UNS_OP5494_3_n_585));
  HAX1 inc_ADD_UNS_OP5494_3_g892(.A (inc_ADD_UNS_OP5494_3_n_591), .B
       (csr_minstret[22]), .S (n_5901), .CO
       (inc_ADD_UNS_OP5494_3_n_588));
  HAX2 inc_ADD_UNS_OP5494_3_g893(.A (inc_ADD_UNS_OP5494_3_n_594), .B
       (csr_minstret[21]), .S (n_5903), .CO
       (inc_ADD_UNS_OP5494_3_n_591));
  NO2I1X1 inc_ADD_UNS_OP5494_3_g895(.B (inc_ADD_UNS_OP5494_3_n_599),
       .AN (csr_minstret[20]), .Q (inc_ADD_UNS_OP5494_3_n_594));
  EO2X0 inc_ADD_UNS_OP5494_3_g897(.A (inc_ADD_UNS_OP5494_3_n_604), .B
       (csr_minstret[19]), .Q (n_5907));
  NA2X1 inc_ADD_UNS_OP5494_3_g898(.A (inc_ADD_UNS_OP5494_3_n_604), .B
       (csr_minstret[19]), .Q (inc_ADD_UNS_OP5494_3_n_599));
  EO2X1 inc_ADD_UNS_OP5494_3_g899(.A (inc_ADD_UNS_OP5494_3_n_607), .B
       (csr_minstret[18]), .Q (n_5909));
  AND4X1 inc_ADD_UNS_OP5494_3_g900(.A (inc_ADD_UNS_OP5494_3_n_613), .B
       (csr_minstret[16]), .C (csr_minstret[17]), .D
       (csr_minstret[18]), .Q (inc_ADD_UNS_OP5494_3_n_604));
  HAX1 inc_ADD_UNS_OP5494_3_g901(.A (inc_ADD_UNS_OP5494_3_n_610), .B
       (csr_minstret[17]), .S (n_5911), .CO
       (inc_ADD_UNS_OP5494_3_n_607));
  HAX1 inc_ADD_UNS_OP5494_3_g902(.A (inc_ADD_UNS_OP5494_3_n_613), .B
       (csr_minstret[16]), .S (n_5913), .CO
       (inc_ADD_UNS_OP5494_3_n_610));
  HAX2 inc_ADD_UNS_OP5494_3_g903(.A (inc_ADD_UNS_OP5494_3_n_616), .B
       (csr_minstret[15]), .S (n_5915), .CO
       (inc_ADD_UNS_OP5494_3_n_613));
  EO2X0 inc_ADD_UNS_OP5494_3_g904(.A (inc_ADD_UNS_OP5494_3_n_736), .B
       (csr_minstret[14]), .Q (n_5917));
  AND2X2 inc_ADD_UNS_OP5494_3_g905(.A (inc_ADD_UNS_OP5494_3_n_736), .B
       (csr_minstret[14]), .Q (inc_ADD_UNS_OP5494_3_n_616));
  EO2X0 inc_ADD_UNS_OP5494_3_g906(.A (inc_ADD_UNS_OP5494_3_n_737), .B
       (csr_minstret[13]), .Q (n_5919));
  EO2X0 inc_ADD_UNS_OP5494_3_g909(.A (inc_ADD_UNS_OP5494_3_n_631), .B
       (csr_minstret[12]), .Q (n_5921));
  NO2I1X1 inc_ADD_UNS_OP5494_3_g913(.B (inc_ADD_UNS_OP5494_3_n_636),
       .AN (csr_minstret[11]), .Q (inc_ADD_UNS_OP5494_3_n_631));
  EO2X0 inc_ADD_UNS_OP5494_3_g915(.A (inc_ADD_UNS_OP5494_3_n_641), .B
       (csr_minstret[10]), .Q (n_5925));
  NA2X2 inc_ADD_UNS_OP5494_3_g916(.A (inc_ADD_UNS_OP5494_3_n_641), .B
       (csr_minstret[10]), .Q (inc_ADD_UNS_OP5494_3_n_636));
  NO2I1X1 inc_ADD_UNS_OP5494_3_g918(.B (inc_ADD_UNS_OP5494_3_n_646),
       .AN (csr_minstret[9]), .Q (inc_ADD_UNS_OP5494_3_n_641));
  EO2X0 inc_ADD_UNS_OP5494_3_g920(.A (inc_ADD_UNS_OP5494_3_n_651), .B
       (csr_minstret[8]), .Q (n_5929));
  NA2X1 inc_ADD_UNS_OP5494_3_g921(.A (inc_ADD_UNS_OP5494_3_n_651), .B
       (csr_minstret[8]), .Q (inc_ADD_UNS_OP5494_3_n_646));
  EO2X0 inc_ADD_UNS_OP5494_3_g922(.A (inc_ADD_UNS_OP5494_3_n_740), .B
       (csr_minstret[7]), .Q (n_5931));
  AND2X1 inc_ADD_UNS_OP5494_3_g923(.A (inc_ADD_UNS_OP5494_3_n_740), .B
       (csr_minstret[7]), .Q (inc_ADD_UNS_OP5494_3_n_651));
  EO2X0 inc_ADD_UNS_OP5494_3_g924(.A (inc_ADD_UNS_OP5494_3_n_661), .B
       (csr_minstret[6]), .Q (n_5933));
  EO2X1 inc_ADD_UNS_OP5494_3_g927(.A (inc_ADD_UNS_OP5494_3_n_664), .B
       (csr_minstret[5]), .Q (n_5935));
  AND5X2 inc_ADD_UNS_OP5494_3_g928(.A (inc_ADD_UNS_OP5494_3_n_673), .B
       (csr_minstret[2]), .C (csr_minstret[3]), .D (csr_minstret[4]),
       .E (csr_minstret[5]), .Q (inc_ADD_UNS_OP5494_3_n_661));
  HAX1 inc_ADD_UNS_OP5494_3_g929(.A (inc_ADD_UNS_OP5494_3_n_667), .B
       (csr_minstret[4]), .S (n_5937), .CO
       (inc_ADD_UNS_OP5494_3_n_664));
  HAX1 inc_ADD_UNS_OP5494_3_g930(.A (inc_ADD_UNS_OP5494_3_n_670), .B
       (csr_minstret[3]), .S (n_5939), .CO
       (inc_ADD_UNS_OP5494_3_n_667));
  HAX1 inc_ADD_UNS_OP5494_3_g931(.A (inc_ADD_UNS_OP5494_3_n_673), .B
       (csr_minstret[2]), .S (n_5941), .CO
       (inc_ADD_UNS_OP5494_3_n_670));
  HAX1 inc_ADD_UNS_OP5494_3_g932(.A (inc_ADD_UNS_OP5494_3_n_676), .B
       (csr_minstret[1]), .S (n_5943), .CO
       (inc_ADD_UNS_OP5494_3_n_673));
  EO2X0 inc_ADD_UNS_OP5494_3_g933(.A (n_6239), .B (csr_minstret[0]), .Q
       (n_5945));
  AND2X2 inc_ADD_UNS_OP5494_3_g934(.A (n_6239), .B (csr_minstret[0]),
       .Q (inc_ADD_UNS_OP5494_3_n_676));
  EO2X1 inc_ADD_UNS_OP5494_3_g2(.A (inc_ADD_UNS_OP5494_3_n_455), .B
       (csr_minstret[62]), .Q (n_5821));
  EN2X0 inc_ADD_UNS_OP5494_3_g937(.A (inc_ADD_UNS_OP5494_3_n_483), .B
       (csr_minstret[50]), .Q (n_5845));
  EN2X0 inc_ADD_UNS_OP5494_3_g938(.A (inc_ADD_UNS_OP5494_3_n_493), .B
       (csr_minstret[48]), .Q (n_5849));
  EN2X0 inc_ADD_UNS_OP5494_3_g939(.A (inc_ADD_UNS_OP5494_3_n_503), .B
       (csr_minstret[46]), .Q (n_5853));
  EN2X0 inc_ADD_UNS_OP5494_3_g940(.A (inc_ADD_UNS_OP5494_3_n_513), .B
       (csr_minstret[44]), .Q (n_5857));
  EN2X0 inc_ADD_UNS_OP5494_3_g941(.A (inc_ADD_UNS_OP5494_3_n_572), .B
       (csr_minstret[27]), .Q (n_5891));
  EN2X1 inc_ADD_UNS_OP5494_3_g942(.A (inc_ADD_UNS_OP5494_3_n_599), .B
       (csr_minstret[20]), .Q (n_5905));
  AND2X1 inc_ADD_UNS_OP5494_3_g943(.A (inc_ADD_UNS_OP5494_3_n_737), .B
       (csr_minstret[13]), .Q (inc_ADD_UNS_OP5494_3_n_736));
  AND2X1 inc_ADD_UNS_OP5494_3_g944(.A (inc_ADD_UNS_OP5494_3_n_631), .B
       (csr_minstret[12]), .Q (inc_ADD_UNS_OP5494_3_n_737));
  EN2X0 inc_ADD_UNS_OP5494_3_g945(.A (inc_ADD_UNS_OP5494_3_n_636), .B
       (csr_minstret[11]), .Q (n_5923));
  EN2X0 inc_ADD_UNS_OP5494_3_g946(.A (inc_ADD_UNS_OP5494_3_n_646), .B
       (csr_minstret[9]), .Q (n_5927));
  AND2X1 inc_ADD_UNS_OP5494_3_g947(.A (inc_ADD_UNS_OP5494_3_n_661), .B
       (csr_minstret[6]), .Q (inc_ADD_UNS_OP5494_3_n_740));
  EN2X1 inc_ADD_UNS_OP5494_3_g948(.A (inc_ADD_UNS_OP5494_3_n_452), .B
       (csr_minstret[63]), .Q (n_5819));
  NO2I1X1 inc_ADD_UNS_OP5494_3_g950(.B (inc_ADD_UNS_OP5494_3_n_483),
       .AN (csr_minstret[50]), .Q (inc_ADD_UNS_OP5494_3_n_478));
  HAX2 inc_ADD_UNS_OP5493_6_g828(.A (inc_ADD_UNS_OP5493_6_n_454), .B
       (n_5729), .S (n_5822), .CO (inc_ADD_UNS_OP5493_6_n_452));
  HAX2 inc_ADD_UNS_OP5493_6_g829(.A (inc_ADD_UNS_OP5493_6_n_456), .B
       (n_5730), .S (n_5824), .CO (inc_ADD_UNS_OP5493_6_n_454));
  HAX2 inc_ADD_UNS_OP5493_6_g830(.A (inc_ADD_UNS_OP5493_6_n_458), .B
       (n_5731), .S (n_5826), .CO (inc_ADD_UNS_OP5493_6_n_456));
  HAX2 inc_ADD_UNS_OP5493_6_g831(.A (inc_ADD_UNS_OP5493_6_n_460), .B
       (n_5732), .S (n_5828), .CO (inc_ADD_UNS_OP5493_6_n_458));
  HAX2 inc_ADD_UNS_OP5493_6_g832(.A (inc_ADD_UNS_OP5493_6_n_462), .B
       (n_5733), .S (n_5830), .CO (inc_ADD_UNS_OP5493_6_n_460));
  HAX2 inc_ADD_UNS_OP5493_6_g833(.A (inc_ADD_UNS_OP5493_6_n_464), .B
       (n_5734), .S (n_5832), .CO (inc_ADD_UNS_OP5493_6_n_462));
  HAX2 inc_ADD_UNS_OP5493_6_g834(.A (inc_ADD_UNS_OP5493_6_n_466), .B
       (n_5735), .S (n_5834), .CO (inc_ADD_UNS_OP5493_6_n_464));
  HAX2 inc_ADD_UNS_OP5493_6_g835(.A (inc_ADD_UNS_OP5493_6_n_468), .B
       (n_5736), .S (n_5836), .CO (inc_ADD_UNS_OP5493_6_n_466));
  HAX2 inc_ADD_UNS_OP5493_6_g836(.A (inc_ADD_UNS_OP5493_6_n_470), .B
       (n_5737), .S (n_5838), .CO (inc_ADD_UNS_OP5493_6_n_468));
  HAX2 inc_ADD_UNS_OP5493_6_g837(.A (inc_ADD_UNS_OP5493_6_n_472), .B
       (n_5738), .S (n_5840), .CO (inc_ADD_UNS_OP5493_6_n_470));
  HAX2 inc_ADD_UNS_OP5493_6_g838(.A (inc_ADD_UNS_OP5493_6_n_474), .B
       (n_5739), .S (n_5842), .CO (inc_ADD_UNS_OP5493_6_n_472));
  NO2I1X1 inc_ADD_UNS_OP5493_6_g840(.B (inc_ADD_UNS_OP5493_6_n_741),
       .AN (n_5740), .Q (inc_ADD_UNS_OP5493_6_n_474));
  EO2X0 inc_ADD_UNS_OP5493_6_g845(.A (inc_ADD_UNS_OP5493_6_n_488), .B
       (n_5742), .Q (n_5848));
  NA2X2 inc_ADD_UNS_OP5493_6_g846(.A (inc_ADD_UNS_OP5493_6_n_488), .B
       (n_5742), .Q (inc_ADD_UNS_OP5493_6_n_483));
  EO2X0 inc_ADD_UNS_OP5493_6_g850(.A (inc_ADD_UNS_OP5493_6_n_498), .B
       (n_4538), .Q (n_5852));
  NA2X2 inc_ADD_UNS_OP5493_6_g851(.A (inc_ADD_UNS_OP5493_6_n_498), .B
       (n_4538), .Q (inc_ADD_UNS_OP5493_6_n_493));
  NO2I1X1 inc_ADD_UNS_OP5493_6_g853(.B (inc_ADD_UNS_OP5493_6_n_503),
       .AN (n_4536), .Q (inc_ADD_UNS_OP5493_6_n_498));
  EO2X1 inc_ADD_UNS_OP5493_6_g855(.A (inc_ADD_UNS_OP5493_6_n_508), .B
       (n_5746), .Q (n_5856));
  NA2X1 inc_ADD_UNS_OP5493_6_g856(.A (inc_ADD_UNS_OP5493_6_n_508), .B
       (n_5746), .Q (inc_ADD_UNS_OP5493_6_n_503));
  EO2X1 inc_ADD_UNS_OP5493_6_g857(.A (inc_ADD_UNS_OP5493_6_n_511), .B
       (n_5747), .Q (n_5858));
  AND6X2 inc_ADD_UNS_OP5493_6_g858(.A (inc_ADD_UNS_OP5493_6_n_525), .B
       (n_5749), .C (n_5748), .D (n_5747), .E (n_5751), .F (n_5750), .Q
       (inc_ADD_UNS_OP5493_6_n_508));
  HAX1 inc_ADD_UNS_OP5493_6_g859(.A (inc_ADD_UNS_OP5493_6_n_514), .B
       (n_5748), .S (n_5860), .CO (inc_ADD_UNS_OP5493_6_n_511));
  HAX1 inc_ADD_UNS_OP5493_6_g860(.A (inc_ADD_UNS_OP5493_6_n_517), .B
       (n_5749), .S (n_5862), .CO (inc_ADD_UNS_OP5493_6_n_514));
  HAX1 inc_ADD_UNS_OP5493_6_g861(.A (inc_ADD_UNS_OP5493_6_n_520), .B
       (n_5750), .S (n_5864), .CO (inc_ADD_UNS_OP5493_6_n_517));
  HAX1 inc_ADD_UNS_OP5493_6_g862(.A (inc_ADD_UNS_OP5493_6_n_525), .B
       (n_5751), .S (n_5866), .CO (inc_ADD_UNS_OP5493_6_n_520));
  EO2X1 inc_ADD_UNS_OP5493_6_g863(.A (inc_ADD_UNS_OP5493_6_n_528), .B
       (n_6726), .Q (n_5868));
  AND5X1 inc_ADD_UNS_OP5493_6_g864(.A (inc_ADD_UNS_OP5493_6_n_537), .B
       (n_4535), .C (n_6730), .D (n_6726), .E (n_6731), .Q
       (inc_ADD_UNS_OP5493_6_n_525));
  HAX1 inc_ADD_UNS_OP5493_6_g865(.A (inc_ADD_UNS_OP5493_6_n_531), .B
       (n_6730), .S (n_5870), .CO (inc_ADD_UNS_OP5493_6_n_528));
  HAX1 inc_ADD_UNS_OP5493_6_g866(.A (inc_ADD_UNS_OP5493_6_n_534), .B
       (n_6731), .S (n_5872), .CO (inc_ADD_UNS_OP5493_6_n_531));
  HAX1 inc_ADD_UNS_OP5493_6_g867(.A (inc_ADD_UNS_OP5493_6_n_537), .B
       (n_4535), .S (n_5874), .CO (inc_ADD_UNS_OP5493_6_n_534));
  HAX1 inc_ADD_UNS_OP5493_6_g868(.A (inc_ADD_UNS_OP5493_6_n_540), .B
       (n_5987), .S (n_5876), .CO (inc_ADD_UNS_OP5493_6_n_537));
  HAX1 inc_ADD_UNS_OP5493_6_g869(.A (inc_ADD_UNS_OP5493_6_n_542), .B
       (n_5988), .S (n_5878), .CO (inc_ADD_UNS_OP5493_6_n_540));
  EO2X1 inc_ADD_UNS_OP5493_6_g870(.A (inc_ADD_UNS_OP5493_6_n_545), .B
       (n_6724), .Q (n_5880));
  AND3X1 inc_ADD_UNS_OP5493_6_g871(.A (inc_ADD_UNS_OP5493_6_n_550), .B
       (n_6724), .C (n_4534), .Q (inc_ADD_UNS_OP5493_6_n_542));
  HAX1 inc_ADD_UNS_OP5493_6_g872(.A (inc_ADD_UNS_OP5493_6_n_550), .B
       (n_4534), .S (n_5882), .CO (inc_ADD_UNS_OP5493_6_n_545));
  EO2X1 inc_ADD_UNS_OP5493_6_g873(.A (inc_ADD_UNS_OP5493_6_n_553), .B
       (csr_minstret[31]), .Q (n_5884));
  AND3X1 inc_ADD_UNS_OP5493_6_g874(.A (inc_ADD_UNS_OP5493_6_n_558), .B
       (csr_minstret[30]), .C (csr_minstret[31]), .Q
       (inc_ADD_UNS_OP5493_6_n_550));
  HAX1 inc_ADD_UNS_OP5493_6_g875(.A (inc_ADD_UNS_OP5493_6_n_558), .B
       (csr_minstret[30]), .S (n_5886), .CO
       (inc_ADD_UNS_OP5493_6_n_553));
  EO2X0 inc_ADD_UNS_OP5493_6_g876(.A (inc_ADD_UNS_OP5493_6_n_563), .B
       (csr_minstret[29]), .Q (n_5888));
  AND2X2 inc_ADD_UNS_OP5493_6_g877(.A (inc_ADD_UNS_OP5493_6_n_563), .B
       (csr_minstret[29]), .Q (inc_ADD_UNS_OP5493_6_n_558));
  EO2X0 inc_ADD_UNS_OP5493_6_g878(.A (inc_ADD_UNS_OP5493_6_n_568), .B
       (csr_minstret[28]), .Q (n_5890));
  AND2X2 inc_ADD_UNS_OP5493_6_g879(.A (inc_ADD_UNS_OP5493_6_n_568), .B
       (csr_minstret[28]), .Q (inc_ADD_UNS_OP5493_6_n_563));
  EO2X1 inc_ADD_UNS_OP5493_6_g880(.A (inc_ADD_UNS_OP5493_6_n_571), .B
       (csr_minstret[27]), .Q (n_5892));
  AND3X1 inc_ADD_UNS_OP5493_6_g881(.A (inc_ADD_UNS_OP5493_6_n_576), .B
       (csr_minstret[26]), .C (csr_minstret[27]), .Q
       (inc_ADD_UNS_OP5493_6_n_568));
  HAX1 inc_ADD_UNS_OP5493_6_g882(.A (inc_ADD_UNS_OP5493_6_n_576), .B
       (csr_minstret[26]), .S (n_5894), .CO
       (inc_ADD_UNS_OP5493_6_n_571));
  EO2X0 inc_ADD_UNS_OP5493_6_g883(.A (inc_ADD_UNS_OP5493_6_n_581), .B
       (csr_minstret[25]), .Q (n_5896));
  AND2X2 inc_ADD_UNS_OP5493_6_g884(.A (inc_ADD_UNS_OP5493_6_n_581), .B
       (csr_minstret[25]), .Q (inc_ADD_UNS_OP5493_6_n_576));
  EO2X0 inc_ADD_UNS_OP5493_6_g885(.A (inc_ADD_UNS_OP5493_6_n_586), .B
       (csr_minstret[24]), .Q (n_5898));
  AND2X2 inc_ADD_UNS_OP5493_6_g886(.A (inc_ADD_UNS_OP5493_6_n_586), .B
       (csr_minstret[24]), .Q (inc_ADD_UNS_OP5493_6_n_581));
  EO2X0 inc_ADD_UNS_OP5493_6_g887(.A (inc_ADD_UNS_OP5493_6_n_591), .B
       (csr_minstret[23]), .Q (n_5900));
  EO2X1 inc_ADD_UNS_OP5493_6_g889(.A (inc_ADD_UNS_OP5493_6_n_594), .B
       (csr_minstret[22]), .Q (n_5902));
  AND3X1 inc_ADD_UNS_OP5493_6_g890(.A (inc_ADD_UNS_OP5493_6_n_599), .B
       (csr_minstret[21]), .C (csr_minstret[22]), .Q
       (inc_ADD_UNS_OP5493_6_n_591));
  HAX1 inc_ADD_UNS_OP5493_6_g891(.A (inc_ADD_UNS_OP5493_6_n_599), .B
       (csr_minstret[21]), .S (n_5904), .CO
       (inc_ADD_UNS_OP5493_6_n_594));
  EO2X1 inc_ADD_UNS_OP5493_6_g892(.A (inc_ADD_UNS_OP5493_6_n_602), .B
       (csr_minstret[20]), .Q (n_5906));
  AND3X1 inc_ADD_UNS_OP5493_6_g893(.A (inc_ADD_UNS_OP5493_6_n_607), .B
       (csr_minstret[19]), .C (csr_minstret[20]), .Q
       (inc_ADD_UNS_OP5493_6_n_599));
  HAX1 inc_ADD_UNS_OP5493_6_g894(.A (inc_ADD_UNS_OP5493_6_n_607), .B
       (csr_minstret[19]), .S (n_5908), .CO
       (inc_ADD_UNS_OP5493_6_n_602));
  EO2X0 inc_ADD_UNS_OP5493_6_g895(.A (inc_ADD_UNS_OP5493_6_n_610), .B
       (csr_minstret[18]), .Q (n_5910));
  AND2X2 inc_ADD_UNS_OP5493_6_g896(.A (inc_ADD_UNS_OP5493_6_n_610), .B
       (csr_minstret[18]), .Q (inc_ADD_UNS_OP5493_6_n_607));
  HAX2 inc_ADD_UNS_OP5493_6_g897(.A (inc_ADD_UNS_OP5493_6_n_613), .B
       (csr_minstret[17]), .S (n_5912), .CO
       (inc_ADD_UNS_OP5493_6_n_610));
  EO2X1 inc_ADD_UNS_OP5493_6_g898(.A (inc_ADD_UNS_OP5493_6_n_616), .B
       (csr_minstret[16]), .Q (n_5914));
  AND4X1 inc_ADD_UNS_OP5493_6_g899(.A (inc_ADD_UNS_OP5493_6_n_622), .B
       (csr_minstret[14]), .C (csr_minstret[15]), .D
       (csr_minstret[16]), .Q (inc_ADD_UNS_OP5493_6_n_613));
  HAX1 inc_ADD_UNS_OP5493_6_g900(.A (inc_ADD_UNS_OP5493_6_n_619), .B
       (csr_minstret[15]), .S (n_5916), .CO
       (inc_ADD_UNS_OP5493_6_n_616));
  HAX1 inc_ADD_UNS_OP5493_6_g901(.A (inc_ADD_UNS_OP5493_6_n_622), .B
       (csr_minstret[14]), .S (n_5918), .CO
       (inc_ADD_UNS_OP5493_6_n_619));
  HAX2 inc_ADD_UNS_OP5493_6_g902(.A (inc_ADD_UNS_OP5493_6_n_625), .B
       (csr_minstret[13]), .S (n_5920), .CO
       (inc_ADD_UNS_OP5493_6_n_622));
  EO2X0 inc_ADD_UNS_OP5493_6_g903(.A (inc_ADD_UNS_OP5493_6_n_630), .B
       (csr_minstret[12]), .Q (n_5922));
  AND2X2 inc_ADD_UNS_OP5493_6_g904(.A (inc_ADD_UNS_OP5493_6_n_630), .B
       (csr_minstret[12]), .Q (inc_ADD_UNS_OP5493_6_n_625));
  NO2I1X1 inc_ADD_UNS_OP5493_6_g906(.B (inc_ADD_UNS_OP5493_6_n_635),
       .AN (csr_minstret[11]), .Q (inc_ADD_UNS_OP5493_6_n_630));
  EO2X0 inc_ADD_UNS_OP5493_6_g908(.A (inc_ADD_UNS_OP5493_6_n_737), .B
       (csr_minstret[10]), .Q (n_5926));
  NA2X1 inc_ADD_UNS_OP5493_6_g909(.A (inc_ADD_UNS_OP5493_6_n_737), .B
       (csr_minstret[10]), .Q (inc_ADD_UNS_OP5493_6_n_635));
  EO2X0 inc_ADD_UNS_OP5493_6_g910(.A (inc_ADD_UNS_OP5493_6_n_738), .B
       (csr_minstret[9]), .Q (n_5928));
  EO2X0 inc_ADD_UNS_OP5493_6_g913(.A (inc_ADD_UNS_OP5493_6_n_650), .B
       (csr_minstret[8]), .Q (n_5930));
  NO2I1X1 inc_ADD_UNS_OP5493_6_g917(.B (inc_ADD_UNS_OP5493_6_n_655),
       .AN (csr_minstret[7]), .Q (inc_ADD_UNS_OP5493_6_n_650));
  EO2X0 inc_ADD_UNS_OP5493_6_g919(.A (inc_ADD_UNS_OP5493_6_n_660), .B
       (csr_minstret[6]), .Q (n_5934));
  NA2X1 inc_ADD_UNS_OP5493_6_g920(.A (inc_ADD_UNS_OP5493_6_n_660), .B
       (csr_minstret[6]), .Q (inc_ADD_UNS_OP5493_6_n_655));
  EO2X0 inc_ADD_UNS_OP5493_6_g921(.A (inc_ADD_UNS_OP5493_6_n_665), .B
       (csr_minstret[5]), .Q (n_5936));
  AND2X2 inc_ADD_UNS_OP5493_6_g922(.A (inc_ADD_UNS_OP5493_6_n_665), .B
       (csr_minstret[5]), .Q (inc_ADD_UNS_OP5493_6_n_660));
  EO2X1 inc_ADD_UNS_OP5493_6_g923(.A (inc_ADD_UNS_OP5493_6_n_668), .B
       (csr_minstret[4]), .Q (n_5938));
  AND6X1 inc_ADD_UNS_OP5493_6_g924(.A (n_6239), .B (csr_minstret[1]),
       .C (csr_minstret[2]), .D (csr_minstret[0]), .E
       (csr_minstret[3]), .F (csr_minstret[4]), .Q
       (inc_ADD_UNS_OP5493_6_n_665));
  HAX1 inc_ADD_UNS_OP5493_6_g925(.A (inc_ADD_UNS_OP5493_6_n_671), .B
       (csr_minstret[3]), .S (n_5940), .CO
       (inc_ADD_UNS_OP5493_6_n_668));
  HAX1 inc_ADD_UNS_OP5493_6_g926(.A (inc_ADD_UNS_OP5493_6_n_674), .B
       (csr_minstret[2]), .S (n_5942), .CO
       (inc_ADD_UNS_OP5493_6_n_671));
  HAX1 inc_ADD_UNS_OP5493_6_g927(.A (inc_ADD_UNS_OP5493_6_n_677), .B
       (csr_minstret[1]), .S (n_5944), .CO
       (inc_ADD_UNS_OP5493_6_n_674));
  HAX1 inc_ADD_UNS_OP5493_6_g928(.A (n_6239), .B (csr_minstret[0]), .S
       (n_5946), .CO (inc_ADD_UNS_OP5493_6_n_677));
  EN2X1 inc_ADD_UNS_OP5493_6_g2(.A (inc_ADD_UNS_OP5493_6_n_741), .B
       (n_5740), .Q (n_5844));
  EN2X0 inc_ADD_UNS_OP5493_6_g931(.A (inc_ADD_UNS_OP5493_6_n_483), .B
       (n_5741), .Q (n_5846));
  EN2X0 inc_ADD_UNS_OP5493_6_g932(.A (inc_ADD_UNS_OP5493_6_n_493), .B
       (n_5743), .Q (n_5850));
  EN2X1 inc_ADD_UNS_OP5493_6_g933(.A (inc_ADD_UNS_OP5493_6_n_503), .B
       (n_4536), .Q (n_5854));
  EN2X0 inc_ADD_UNS_OP5493_6_g934(.A (inc_ADD_UNS_OP5493_6_n_635), .B
       (csr_minstret[11]), .Q (n_5924));
  AND2X1 inc_ADD_UNS_OP5493_6_g935(.A (inc_ADD_UNS_OP5493_6_n_738), .B
       (csr_minstret[9]), .Q (inc_ADD_UNS_OP5493_6_n_737));
  AND2X1 inc_ADD_UNS_OP5493_6_g936(.A (inc_ADD_UNS_OP5493_6_n_650), .B
       (csr_minstret[8]), .Q (inc_ADD_UNS_OP5493_6_n_738));
  EN2X0 inc_ADD_UNS_OP5493_6_g937(.A (inc_ADD_UNS_OP5493_6_n_655), .B
       (csr_minstret[7]), .Q (n_5932));
  EO2X1 inc_ADD_UNS_OP5493_6_g938(.A (inc_ADD_UNS_OP5493_6_n_452), .B
       (n_5985), .Q (n_5820));
  NA2I1X2 inc_ADD_UNS_OP5493_6_g939(.B (n_5741), .AN
       (inc_ADD_UNS_OP5493_6_n_483), .Q (inc_ADD_UNS_OP5493_6_n_741));
  NO2I1X2 inc_ADD_UNS_OP5493_6_g941(.B (inc_ADD_UNS_OP5493_6_n_493),
       .AN (n_5743), .Q (inc_ADD_UNS_OP5493_6_n_488));
  AND2X1 inc_ADD_UNS_OP5493_6_g943(.A (inc_ADD_UNS_OP5493_6_n_591), .B
       (csr_minstret[23]), .Q (inc_ADD_UNS_OP5493_6_n_586));
  EO2X1 add_1545_30_g1211(.A (add_1545_30_n_700), .B (csr_mtvec[27]),
       .Q (n_6189));
  EO2X1 add_1545_30_g1212(.A (add_1545_30_n_703), .B (csr_mtvec[23]),
       .Q (n_6193));
  HAX1 add_1545_30_g1213(.A (add_1545_30_n_710), .B (csr_mtvec[26]), .S
       (n_6190), .CO (add_1545_30_n_700));
  EO2X1 add_1545_30_g1214(.A (add_1545_30_n_706), .B (csr_mtvec[19]),
       .Q (n_6197));
  HAX1 add_1545_30_g1215(.A (add_1545_30_n_719), .B (csr_mtvec[22]), .S
       (n_6194), .CO (add_1545_30_n_703));
  EO2X1 add_1545_30_g1216(.A (add_1545_30_n_712), .B (csr_mtvec[15]),
       .Q (n_6201));
  HAX1 add_1545_30_g1217(.A (add_1545_30_n_721), .B (csr_mtvec[18]), .S
       (n_6198), .CO (add_1545_30_n_706));
  EO2X1 add_1545_30_g1218(.A (add_1545_30_n_715), .B (csr_mtvec[31]),
       .Q (n_6185));
  EO2X1 add_1545_30_g1219(.A (add_1545_30_n_717), .B (csr_mtvec[11]),
       .Q (n_6205));
  HAX1 add_1545_30_g1220(.A (add_1545_30_n_725), .B (csr_mtvec[25]), .S
       (n_6191), .CO (add_1545_30_n_710));
  HAX1 add_1545_30_g1221(.A (add_1545_30_n_727), .B (csr_mtvec[14]), .S
       (n_6202), .CO (add_1545_30_n_712));
  EO2X1 add_1545_30_g1222(.A (add_1545_30_n_723), .B (csr_mtvec[29]),
       .Q (n_6187));
  HAX1 add_1545_30_g1223(.A (add_1545_30_n_732), .B (csr_mtvec[30]), .S
       (n_6186), .CO (add_1545_30_n_715));
  HAX1 add_1545_30_g1224(.A (add_1545_30_n_729), .B (csr_mtvec[10]), .S
       (n_6206), .CO (add_1545_30_n_717));
  HAX1 add_1545_30_g1225(.A (add_1545_30_n_731), .B (csr_mtvec[21]), .S
       (n_6195), .CO (add_1545_30_n_719));
  HAX1 add_1545_30_g1226(.A (add_1545_30_n_737), .B (csr_mtvec[17]), .S
       (n_6199), .CO (add_1545_30_n_721));
  HAX1 add_1545_30_g1227(.A (add_1545_30_n_738), .B (csr_mtvec[28]), .S
       (n_6188), .CO (add_1545_30_n_723));
  HAX1 add_1545_30_g1228(.A (add_1545_30_n_746), .B (csr_mtvec[24]), .S
       (n_6192), .CO (add_1545_30_n_725));
  HAX1 add_1545_30_g1229(.A (add_1545_30_n_745), .B (csr_mtvec[13]), .S
       (n_6203), .CO (add_1545_30_n_727));
  HAX1 add_1545_30_g1230(.A (add_1545_30_n_753), .B (csr_mtvec[9]), .S
       (n_6207), .CO (add_1545_30_n_729));
  HAX1 add_1545_30_g1231(.A (add_1545_30_n_754), .B (csr_mtvec[20]), .S
       (n_6196), .CO (add_1545_30_n_731));
  AND3X1 add_1545_30_g1232(.A (add_1545_30_n_738), .B (csr_mtvec[28]),
       .C (csr_mtvec[29]), .Q (add_1545_30_n_732));
  HAX1 add_1545_30_g1233(.A (add_1545_30_n_760), .B (csr_mtvec[16]), .S
       (n_6200), .CO (add_1545_30_n_737));
  AND5X1 add_1545_30_g1234(.A (add_1545_30_n_746), .B (csr_mtvec[24]),
       .C (csr_mtvec[25]), .D (csr_mtvec[27]), .E (csr_mtvec[26]), .Q
       (add_1545_30_n_738));
  HAX1 add_1545_30_g1235(.A (add_1545_30_n_766), .B (csr_mtvec[12]), .S
       (n_6204), .CO (add_1545_30_n_745));
  AND5X1 add_1545_30_g1236(.A (add_1545_30_n_754), .B (csr_mtvec[20]),
       .C (csr_mtvec[21]), .D (csr_mtvec[23]), .E (csr_mtvec[22]), .Q
       (add_1545_30_n_746));
  HAX1 add_1545_30_g1237(.A (add_1545_30_n_772), .B (csr_mtvec[8]), .S
       (n_6208), .CO (add_1545_30_n_753));
  AND5X1 add_1545_30_g1238(.A (add_1545_30_n_760), .B (csr_mtvec[16]),
       .C (csr_mtvec[17]), .D (csr_mtvec[19]), .E (csr_mtvec[18]), .Q
       (add_1545_30_n_754));
  AND5X1 add_1545_30_g1239(.A (add_1545_30_n_766), .B (csr_mtvec[12]),
       .C (csr_mtvec[13]), .D (csr_mtvec[15]), .E (csr_mtvec[14]), .Q
       (add_1545_30_n_760));
  AND5X1 add_1545_30_g1240(.A (add_1545_30_n_772), .B (csr_mtvec[8]),
       .C (csr_mtvec[9]), .D (csr_mtvec[11]), .E (csr_mtvec[10]), .Q
       (add_1545_30_n_766));
  HAX1 add_1545_30_g1241(.A (add_1545_30_n_775), .B (csr_mtvec[7]), .S
       (n_6209), .CO (add_1545_30_n_772));
  FAX0 add_1545_30_g1242(.A (add_1545_30_n_777), .B
       (csr_mcause_code[4]), .CI (csr_mtvec[6]), .S (n_6210), .CO
       (add_1545_30_n_775));
  FAX1 add_1545_30_g1243(.A (csr_mtvec[5]), .B (csr_mcause_code[3]),
       .CI (add_1545_30_n_779), .S (n_6211), .CO (add_1545_30_n_777));
  FAX1 add_1545_30_g1244(.A (csr_mtvec[4]), .B (csr_mcause_code[2]),
       .CI (add_1545_30_n_781), .S (n_6212), .CO (add_1545_30_n_779));
  FAX1 add_1545_30_g1245(.A (csr_mtvec[3]), .B (csr_mcause_code[1]),
       .CI (add_1545_30_n_783), .S (n_6213), .CO (add_1545_30_n_781));
  HAX1 add_1545_30_g1246(.A (csr_mcause_code[0]), .B (csr_mtvec[2]), .S
       (n_6214), .CO (add_1545_30_n_783));
  EO2X1 add_459_21_g1199(.A (add_459_21_n_755), .B
       (program_counter[31]), .Q (n_5603));
  EO2X1 add_459_21_g1200(.A (add_459_21_n_758), .B
       (program_counter[27]), .Q (n_5599));
  HAX1 add_459_21_g1201(.A (add_459_21_n_764), .B
       (program_counter[30]), .S (n_5602), .CO (add_459_21_n_755));
  EO2X1 add_459_21_g1202(.A (add_459_21_n_761), .B
       (program_counter[23]), .Q (n_5595));
  HAX1 add_459_21_g1203(.A (add_459_21_n_771), .B
       (program_counter[26]), .S (n_5598), .CO (add_459_21_n_758));
  EO2X1 add_459_21_g1204(.A (add_459_21_n_766), .B
       (program_counter[19]), .Q (n_5591));
  HAX1 add_459_21_g1205(.A (add_459_21_n_774), .B
       (program_counter[22]), .S (n_5594), .CO (add_459_21_n_761));
  EO2X1 add_459_21_g1206(.A (add_459_21_n_769), .B
       (program_counter[15]), .Q (n_5587));
  HAX1 add_459_21_g1207(.A (add_459_21_n_782), .B
       (program_counter[29]), .S (n_5601), .CO (add_459_21_n_764));
  HAX1 add_459_21_g1208(.A (add_459_21_n_780), .B
       (program_counter[18]), .S (n_5590), .CO (add_459_21_n_766));
  EO2X1 add_459_21_g1209(.A (add_459_21_n_776), .B
       (program_counter[11]), .Q (n_5583));
  HAX1 add_459_21_g1210(.A (add_459_21_n_786), .B
       (program_counter[14]), .S (n_5586), .CO (add_459_21_n_769));
  HAX1 add_459_21_g1211(.A (add_459_21_n_784), .B
       (program_counter[25]), .S (n_5597), .CO (add_459_21_n_771));
  EO2X1 add_459_21_g1212(.A (add_459_21_n_778), .B
       (program_counter[7]), .Q (n_5579));
  HAX1 add_459_21_g1213(.A (add_459_21_n_790), .B
       (program_counter[21]), .S (n_5593), .CO (add_459_21_n_774));
  HAX1 add_459_21_g1214(.A (add_459_21_n_788), .B
       (program_counter[10]), .S (n_5582), .CO (add_459_21_n_776));
  HAX1 add_459_21_g1215(.A (add_459_21_n_792), .B (program_counter[6]),
       .S (n_5578), .CO (add_459_21_n_778));
  HAX1 add_459_21_g1216(.A (add_459_21_n_794), .B
       (program_counter[17]), .S (n_5589), .CO (add_459_21_n_780));
  HAX1 add_459_21_g1217(.A (add_459_21_n_795), .B
       (program_counter[28]), .S (n_5600), .CO (add_459_21_n_782));
  HAX1 add_459_21_g1218(.A (add_459_21_n_803), .B
       (program_counter[24]), .S (n_5596), .CO (add_459_21_n_784));
  HAX1 add_459_21_g1219(.A (add_459_21_n_802), .B
       (program_counter[13]), .S (n_5585), .CO (add_459_21_n_786));
  HAX1 add_459_21_g1220(.A (add_459_21_n_810), .B (program_counter[9]),
       .S (n_5581), .CO (add_459_21_n_788));
  HAX1 add_459_21_g1221(.A (add_459_21_n_811), .B
       (program_counter[20]), .S (n_5592), .CO (add_459_21_n_790));
  HAX1 add_459_21_g1222(.A (add_459_21_n_818), .B (program_counter[5]),
       .S (n_5577), .CO (add_459_21_n_792));
  HAX1 add_459_21_g1223(.A (add_459_21_n_819), .B
       (program_counter[16]), .S (n_5588), .CO (add_459_21_n_794));
  AND5X1 add_459_21_g1224(.A (add_459_21_n_803), .B
       (program_counter[24]), .C (program_counter[25]), .D
       (program_counter[27]), .E (program_counter[26]), .Q
       (add_459_21_n_795));
  HAX1 add_459_21_g1225(.A (add_459_21_n_825), .B
       (program_counter[12]), .S (n_5584), .CO (add_459_21_n_802));
  AND5X1 add_459_21_g1226(.A (add_459_21_n_811), .B
       (program_counter[20]), .C (program_counter[21]), .D
       (program_counter[23]), .E (program_counter[22]), .Q
       (add_459_21_n_803));
  HAX1 add_459_21_g1227(.A (add_459_21_n_831), .B (program_counter[8]),
       .S (n_5580), .CO (add_459_21_n_810));
  AND5X1 add_459_21_g1228(.A (add_459_21_n_819), .B
       (program_counter[16]), .C (program_counter[17]), .D
       (program_counter[19]), .E (program_counter[18]), .Q
       (add_459_21_n_811));
  HAX1 add_459_21_g1229(.A (add_459_21_n_837), .B (program_counter[4]),
       .S (n_5576), .CO (add_459_21_n_818));
  AND5X1 add_459_21_g1230(.A (add_459_21_n_825), .B
       (program_counter[12]), .C (program_counter[13]), .D
       (program_counter[15]), .E (program_counter[14]), .Q
       (add_459_21_n_819));
  AND5X1 add_459_21_g1231(.A (add_459_21_n_831), .B
       (program_counter[8]), .C (program_counter[9]), .D
       (program_counter[11]), .E (program_counter[10]), .Q
       (add_459_21_n_825));
  AND5X1 add_459_21_g1232(.A (add_459_21_n_837), .B
       (program_counter[4]), .C (program_counter[5]), .D
       (program_counter[7]), .E (program_counter[6]), .Q
       (add_459_21_n_831));
  HAX1 add_459_21_g1233(.A (program_counter[2]), .B
       (program_counter[3]), .S (n_5575), .CO (add_459_21_n_837));
  EN2X1 g64021(.A (n_3138), .B (alu_operation_code_39061), .Q (n_6607));
  AO22X1 g64022(.A (n_6453), .B (csr_data_out[5]), .C (n_5577), .D
       (n_4532), .Q (n_6608));
  AN22X1 g64023(.A (n_5574), .B (n_4532), .C (csr_data_out[2]), .D
       (n_6453), .Q (n_6609));
  AN22X1 g64024(.A (n_5575), .B (n_4532), .C (csr_data_out[3]), .D
       (n_6453), .Q (n_6610));
  AN22X1 g64025(.A (program_counter[1]), .B (n_4532), .C
       (csr_data_out[1]), .D (n_6453), .Q (n_6611));
  AN22X1 g64026(.A (n_5583), .B (n_4532), .C (csr_data_out[11]), .D
       (n_6453), .Q (n_6612));
  AO22X1 g64027(.A (n_6453), .B (csr_data_out[7]), .C (n_5579), .D
       (n_4532), .Q (n_6613));
  AO22X1 g64028(.A (n_6453), .B (csr_data_out[8]), .C (n_5580), .D
       (n_4532), .Q (n_6614));
  AO22X1 g64029(.A (n_6453), .B (csr_data_out[10]), .C (n_5582), .D
       (n_4532), .Q (n_6615));
  AN22X1 g64030(.A (n_5581), .B (n_4532), .C (csr_data_out[9]), .D
       (n_6453), .Q (n_6616));
  AO22X1 g64031(.A (n_6453), .B (csr_data_out[4]), .C (n_5576), .D
       (n_4532), .Q (n_6617));
  AO22X1 g64032(.A (n_6453), .B (csr_data_out[6]), .C (n_5578), .D
       (n_4532), .Q (n_6618));
  NA2X1 g64033(.A (csr_data_out[0]), .B (n_6453), .Q (n_6619));
  AN21X1 g64034(.A (n_5723), .B (n_298), .C (n_559), .Q (n_6620));
  AN21X1 g64035(.A (add_463_14_n_900), .B (n_6621), .C
       (add_463_14_n_882), .Q (n_6622));
  AO21X1 g3(.A (add_463_14_n_890), .B (add_463_14_n_696), .C
       (add_463_14_n_893), .Q (n_6621));
  NA2I1X2 g64036(.B (n_3494), .AN (jal_type), .Q (n_6623));
  NO2I1X4 g64037(.B (n_1856), .AN (n_1570), .Q (n_6624));
  NO2I1X4 g64038(.B (n_1851), .AN (n_1570), .Q (n_6625));
  NA5I1X2 g64040(.B (n_4415), .C (n_4391), .D (n_6689), .E (n_6679),
       .AN (n_6636), .Q (n_6627));
  NA6I1X4 g64041(.B (n_3310), .C (n_3309), .D (n_4426), .E (n_3829), .F
       (n_3830), .AN (n_4223), .Q (n_6628));
  NA6I1X4 g64042(.B (n_4367), .C (n_4366), .D (n_6712), .E (n_3797), .F
       (n_3798), .AN (n_4361), .Q (n_6629));
  AND5X1 g64043(.A (n_6657), .B (n_6655), .C (n_3326), .D (n_4196), .E
       (n_3996), .Q (n_6630));
  AND5X1 g64044(.A (n_6658), .B (n_4333), .C (n_3325), .D (n_3972), .E
       (n_3988), .Q (n_6631));
  NA3X1 g64047(.A (n_6678), .B (n_3957), .C (n_3917), .Q (n_6634));
  NA3X1 g64048(.A (n_3914), .B (n_3954), .C (n_3321), .Q (n_6635));
  NA3I2X2 g64049(.C (n_3318), .AN (n_3949), .BN (n_3909), .Q (n_6636));
  NA3X1 g64050(.A (n_3910), .B (n_3950), .C (n_6688), .Q (n_6637));
  NA3X1 g64051(.A (n_3853), .B (n_3854), .C (n_4227), .Q (n_6638));
  NA3X1 g64052(.A (n_3851), .B (n_3852), .C (n_6708), .Q (n_6639));
  NA3X1 g64053(.A (n_3837), .B (n_3855), .C (n_6703), .Q (n_6640));
  NA3X1 g64054(.A (n_3826), .B (n_3834), .C (n_6781), .Q (n_6641));
  AN221X1 g64055(.A (n_6768), .B (n_5288), .C (n_6767), .D (n_5289), .E
       (n_3899), .Q (n_6642));
  AN221X1 g64056(.A (n_3510), .B (n_5299), .C (n_3508), .D (n_5300), .E
       (n_4157), .Q (n_6643));
  AN221X1 g64057(.A (n_3301), .B (n_5171), .C (n_3512), .D (n_5172), .E
       (n_4174), .Q (n_6644));
  AN221X1 g64058(.A (n_3524), .B (n_5332), .C (n_3514), .D (n_5333), .E
       (n_4183), .Q (n_6645));
  AN221X1 g64059(.A (n_3524), .B (n_5301), .C (n_3514), .D (n_5302), .E
       (n_4181), .Q (n_6646));
  AN221X1 g64060(.A (n_3510), .B (n_5330), .C (n_3526), .D (n_5329), .E
       (n_4159), .Q (n_6647));
  AN221X1 g64061(.A (n_3524), .B (n_4712), .C (n_3514), .D (n_4713), .E
       (n_4169), .Q (n_6648));
  AN221X1 g64062(.A (n_3301), .B (n_5450), .C (n_3512), .D (n_5451), .E
       (n_4127), .Q (n_6649));
  AN221X1 g64063(.A (n_3524), .B (n_4619), .C (n_3514), .D (n_4620), .E
       (n_4166), .Q (n_6650));
  AN221X1 g64064(.A (n_3301), .B (n_4830), .C (n_3512), .D (n_4831), .E
       (n_4104), .Q (n_6651));
  AN221X1 g64065(.A (n_3524), .B (n_5084), .C (n_3514), .D (n_5085), .E
       (n_4135), .Q (n_6652));
  AN221X1 g64066(.A (n_3524), .B (n_5518), .C (n_3514), .D (n_5519), .E
       (n_4132), .Q (n_6653));
  AN221X1 g64067(.A (n_3524), .B (n_5363), .C (n_3514), .D (n_5364), .E
       (n_4131), .Q (n_6654));
  AN221X1 g64068(.A (n_3509), .B (n_4835), .C (n_3305), .D (n_4840), .E
       (n_4101), .Q (n_6655));
  AN221X1 g64069(.A (n_3510), .B (n_5082), .C (n_3526), .D (n_5081), .E
       (n_4098), .Q (n_6656));
  AN221X1 g64070(.A (n_3522), .B (n_4842), .C (n_3298), .D (n_4841), .E
       (n_4133), .Q (n_6657));
  AN221X1 g64071(.A (n_3509), .B (n_5517), .C (n_3305), .D (n_5522), .E
       (n_4129), .Q (n_6658));
  AN221X1 g64072(.A (n_3542), .B (n_5313), .C (n_3544), .D (n_5314), .E
       (n_4106), .Q (n_6659));
  AN221X1 g64073(.A (n_3542), .B (n_5344), .C (n_3544), .D (n_5345), .E
       (n_4110), .Q (n_6660));
  AN221X1 g64074(.A (n_3546), .B (n_4733), .C (n_3536), .D (n_4732), .E
       (n_4047), .Q (n_6661));
  AN221X1 g64075(.A (n_3542), .B (n_4724), .C (n_3544), .D (n_4725), .E
       (n_4042), .Q (n_6662));
  AN211X1 g64076(.A (n_3505), .B (n_5046), .C (n_4028), .D (n_3683), .Q
       (n_6663));
  AN221X1 g64077(.A (n_3522), .B (n_5493), .C (n_3298), .D (n_5492), .E
       (n_4025), .Q (n_6664));
  AN221X1 g64078(.A (n_3301), .B (n_4954), .C (n_3512), .D (n_4955), .E
       (n_4018), .Q (n_6665));
  AN221X1 g64079(.A (n_3522), .B (n_4966), .C (n_3298), .D (n_4965), .E
       (n_4017), .Q (n_6666));
  AN221X1 g64080(.A (n_3544), .B (n_5066), .C (n_3542), .D (n_5065), .E
       (n_3960), .Q (n_6667));
  AN221X1 g64081(.A (n_3538), .B (n_5253), .C (n_3540), .D (n_5254), .E
       (n_3937), .Q (n_6668));
  AN221X1 g64082(.A (n_3504), .B (n_5262), .C (n_3547), .D (n_5261), .E
       (n_3935), .Q (n_6669));
  AN221X1 g64083(.A (n_3547), .B (n_5230), .C (n_3504), .D (n_5231), .E
       (n_3930), .Q (n_6670));
  AN221X1 g64084(.A (n_3551), .B (n_5155), .C (n_3549), .D (n_5154), .E
       (n_3968), .Q (n_6671));
  AN221X1 g64085(.A (n_3548), .B (n_5162), .C (n_3557), .D (n_5163), .E
       (n_3967), .Q (n_6672));
  AN221X1 g64086(.A (n_6768), .B (n_5164), .C (n_6767), .D (n_5165), .E
       (n_3966), .Q (n_6673));
  AN221X1 g64087(.A (n_3557), .B (n_5070), .C (n_3548), .D (n_5069), .E
       (n_3963), .Q (n_6674));
  AN221X1 g64088(.A (n_3551), .B (n_5496), .C (n_3549), .D (n_5495), .E
       (n_3962), .Q (n_6675));
  AN221X1 g64089(.A (n_3549), .B (n_5061), .C (n_3551), .D (n_5062), .E
       (n_3920), .Q (n_6676));
  AN221X1 g64090(.A (n_3557), .B (n_5504), .C (n_3548), .D (n_5503), .E
       (n_3958), .Q (n_6677));
  AN221X1 g64091(.A (n_3554), .B (n_5002), .C (n_3553), .D (n_5001), .E
       (n_3956), .Q (n_6678));
  AN221X1 g64092(.A (n_3557), .B (n_4915), .C (n_3548), .D (n_4914), .E
       (n_3946), .Q (n_6679));
  AN221X1 g64093(.A (n_3544), .B (n_5283), .C (n_3542), .D (n_5282), .E
       (n_3901), .Q (n_6680));
  AN221X1 g64094(.A (n_6767), .B (n_5258), .C (n_6768), .D (n_5257), .E
       (n_3895), .Q (n_6681));
  AN221X1 g64095(.A (n_3542), .B (n_5220), .C (n_3544), .D (n_5221), .E
       (n_3893), .Q (n_6682));
  AN221X1 g64096(.A (n_3553), .B (n_5218), .C (n_3554), .D (n_5219), .E
       (n_3932), .Q (n_6683));
  AN221X1 g64097(.A (n_6767), .B (n_5227), .C (n_6768), .D (n_5226), .E
       (n_3971), .Q (n_6684));
  AN221X1 g64098(.A (n_3542), .B (n_5499), .C (n_3544), .D (n_5500), .E
       (n_3923), .Q (n_6685));
  AN221X1 g64099(.A (n_6767), .B (n_5072), .C (n_6768), .D (n_5071), .E
       (n_3965), .Q (n_6686));
  AN221X1 g64100(.A (n_3536), .B (n_5507), .C (n_3546), .D (n_5508), .E
       (n_3919), .Q (n_6687));
  AN221X1 g64101(.A (n_3542), .B (n_4972), .C (n_3544), .D (n_4973), .E
       (n_3911), .Q (n_6688));
  AN221X1 g64102(.A (n_3536), .B (n_4918), .C (n_3546), .D (n_4919), .E
       (n_3907), .Q (n_6689));
  AN221X1 g64103(.A (n_3303), .B (n_4561), .C (n_3526), .D (n_4554), .E
       (n_3886), .Q (n_6690));
  AN221X1 g64104(.A (n_3303), .B (n_4685), .C (n_3505), .D (n_4674), .E
       (n_3875), .Q (n_6691));
  AN221X1 g64105(.A (n_3303), .B (n_4654), .C (n_3505), .D (n_4643), .E
       (n_3868), .Q (n_6692));
  AN221X1 g64106(.A (n_3522), .B (n_4563), .C (n_3505), .D (n_4550), .E
       (n_3888), .Q (n_6693));
  AN221X1 g64107(.A (n_3522), .B (n_4687), .C (n_3507), .D (n_4686), .E
       (n_3874), .Q (n_6694));
  AN221X1 g64108(.A (n_3522), .B (n_4656), .C (n_3507), .D (n_4655), .E
       (n_3869), .Q (n_6695));
  AN221X1 g64109(.A (n_3522), .B (n_4935), .C (n_3507), .D (n_4934), .E
       (n_3881), .Q (n_6696));
  AN222X1 g64110(.A (n_3520), .B (n_5080), .C (n_3518), .D (n_5086), .E
       (n_3517), .F (n_5087), .Q (n_6697));
  AO222X1 g64111(.A (n_3518), .B (n_5489), .C (n_3517), .D (n_5490), .E
       (n_3520), .F (n_5483), .Q (n_6698));
  AO222X1 g64112(.A (n_3518), .B (n_5055), .C (n_3517), .D (n_5056), .E
       (n_3520), .F (n_5049), .Q (n_6699));
  AN221X1 g64113(.A (n_3538), .B (n_4571), .C (n_3540), .D (n_4572), .E
       (n_3866), .Q (n_6700));
  AN221X1 g64114(.A (n_3536), .B (n_4577), .C (n_3546), .D (n_4578), .E
       (n_3863), .Q (n_6701));
  AN221X1 g64115(.A (n_3538), .B (n_4695), .C (n_3540), .D (n_4696), .E
       (n_3858), .Q (n_6702));
  AN221X1 g64116(.A (n_3536), .B (n_4701), .C (n_3546), .D (n_4702), .E
       (n_3838), .Q (n_6703));
  AN221X1 g64117(.A (n_3553), .B (n_4567), .C (n_3554), .D (n_4568), .E
       (n_3850), .Q (n_6704));
  AN221X1 g64118(.A (n_3548), .B (n_4573), .C (n_3557), .D (n_4574), .E
       (n_3841), .Q (n_6705));
  ON221X1 g64119(.A (n_3550), .B (n_3372), .C (n_3552), .D (n_3361), .E
       (n_3847), .Q (n_6706));
  AN221X1 g64120(.A (n_3549), .B (n_4689), .C (n_3551), .D (n_4690), .E
       (n_3845), .Q (n_6707));
  AN221X1 g64121(.A (n_6768), .B (n_4668), .C (n_6767), .D (n_4669), .E
       (n_3836), .Q (n_6708));
  AN211X1 g64123(.A (n_3518), .B (n_4652), .C (n_3592), .D (n_3599), .Q
       (n_6710));
  AN221X1 g64124(.A (n_3549), .B (n_4875), .C (n_3551), .D (n_4876), .E
       (n_3802), .Q (n_6711));
  AN221X1 g64125(.A (n_3536), .B (n_4794), .C (n_3546), .D (n_4795), .E
       (n_3784), .Q (n_6712));
  AN221X1 g64126(.A (n_3553), .B (n_4877), .C (n_3554), .D (n_4878), .E
       (n_6715), .Q (n_6713));
  AN221X1 g64127(.A (n_3553), .B (n_5249), .C (n_3554), .D (n_5250), .E
       (n_3897), .Q (n_6714));
  AO22X2 g64128(.A (n_3542), .B (n_4879), .C (n_3544), .D (n_4880), .Q
       (n_6715));
  AO222X2 g64129(.A (n_6623), .B (instruction[21]), .C (n_3464), .D
       (\instruction[8]_40015 ), .E (n_6453), .F (instruction[16]), .Q
       (n_6716));
  AO222X2 g64130(.A (n_6623), .B (instruction[24]), .C (n_3464), .D
       (\instruction[11]_40800 ), .E (n_6453), .F (instruction[19]), .Q
       (n_6717));
  AO221X2 g64131(.A (n_3394), .B (read_data[1]), .C (n_3393), .D
       (prev_instruction[1]), .E (flush_37507), .Q (n_6718));
  AO22X2 g64132(.A (n_3287), .B (read_data[31]), .C (n_3285), .D
       (prev_instruction[31]), .Q (n_6719));
  AO22X2 g64133(.A (n_3285), .B (prev_instruction[12]), .C (n_3287), .D
       (read_data[12]), .Q (n_6720));
  AO21X2 g64134(.A (n_3285), .B (prev_instruction[13]), .C (n_3409), .Q
       (n_6721));
  AO22X2 g64135(.A (n_3287), .B (read_data[30]), .C (n_3285), .D
       (prev_instruction[30]), .Q (n_6722));
  AO21X4 g64136(.A (n_3392), .B (prev_instruction[20]), .C (n_3396), .Q
       (n_6723));
  AO22X4 g64137(.A (n_1901), .B (csr_data_out[1]), .C (n_1773), .D
       (n_1767), .Q (n_6724));
  NO3I1X1 g64138(.B (n_3140), .C (n_3158), .AN (n_3133), .Q (n_6725));
  AO22X1 g64139(.A (n_1879), .B (csr_data_out[7]), .C
       (\rs1_data[7]_39386 ), .D (n_1586), .Q (n_6726));
  NO5I2X4 g64142(.C (n_3003), .D (n_2819), .E (n_2820), .AN (n_1609),
       .BN (n_1606), .Q (n_6729));
  AO22X2 g64143(.A (n_1899), .B (csr_data_out[6]), .C (n_4466), .D
       (n_1586), .Q (n_6730));
  AO22X2 g64144(.A (n_1873), .B (csr_data_out[5]), .C (n_4461), .D
       (n_1586), .Q (n_6731));
  NA3X1 g64146(.A (n_2396), .B (n_2395), .C (n_6751), .Q (n_6733));
  AN221X1 g64147(.A (n_2196), .B (n_5160), .C (n_2195), .D (n_5159), .E
       (n_2558), .Q (n_6734));
  AN221X1 g64148(.A (n_2181), .B (n_5216), .C (n_2177), .D (n_5217), .E
       (n_2560), .Q (n_6735));
  AN221X1 g64149(.A (n_2196), .B (n_5222), .C (n_2179), .D (n_5218), .E
       (n_2561), .Q (n_6736));
  AO222X1 g64150(.A (n_2159), .B (n_4716), .C (n_1595), .D (n_4708), .E
       (n_2188), .F (n_4705), .Q (n_6737));
  AN221X1 g64151(.A (n_1595), .B (n_4646), .C (n_2188), .D (n_4643), .E
       (n_2719), .Q (n_6738));
  AN221X1 g64152(.A (n_2154), .B (n_5184), .C (n_2156), .D (n_5183), .E
       (n_2786), .Q (n_6739));
  ON221X1 g64153(.A (n_2158), .B (n_1684), .C (n_1597), .D (n_1712), .E
       (n_2351), .Q (n_6740));
  ON221X1 g64154(.A (n_2155), .B (n_1669), .C (n_2157), .D (n_1671), .E
       (n_2571), .Q (n_6741));
  AN221X1 g64155(.A (n_2173), .B (n_5075), .C (n_1600), .D (n_5074), .E
       (n_2503), .Q (n_6742));
  AO222X1 g64156(.A (n_2159), .B (n_4685), .C (n_2160), .D (n_4681), .E
       (n_2164), .F (n_4686), .Q (n_6743));
  AN221X1 g64157(.A (n_2200), .B (n_5021), .C (n_2153), .D (n_5023), .E
       (n_2534), .Q (n_6744));
  AN221X1 g64158(.A (n_2160), .B (n_5270), .C (n_2159), .D (n_5274), .E
       (n_2364), .Q (n_6745));
  AN221X1 g64159(.A (n_2152), .B (n_4962), .C (n_2150), .D (n_4963), .E
       (n_2526), .Q (n_6746));
  AO222X2 g64160(.A (n_2159), .B (n_4809), .C (n_2161), .D (n_4805), .E
       (n_2164), .F (n_4810), .Q (n_6747));
  AN221X1 g64161(.A (n_2181), .B (n_5154), .C (n_2177), .D (n_5155), .E
       (n_2557), .Q (n_6748));
  ON221X1 g64162(.A (n_2158), .B (n_1679), .C (n_1597), .D (n_1713), .E
       (n_2350), .Q (n_6749));
  ON211X1 g64163(.A (n_1601), .B (n_1667), .C (n_2511), .D (n_1858), .Q
       (n_6750));
  AN221X1 g64164(.A (n_2173), .B (n_4765), .C (n_1598), .D (n_4764), .E
       (n_2385), .Q (n_6751));
  AN221X1 g64165(.A (n_2154), .B (n_4781), .C (n_2156), .D (n_4780), .E
       (n_2433), .Q (n_6752));
  AN21X1 g64166(.A (n_1813), .B (n_4797), .C (n_2288), .Q (n_6753));
  AN222X1 g64167(.A (n_2159), .B (n_4747), .C (n_2161), .D (n_4743), .E
       (n_2164), .F (n_4748), .Q (n_6754));
  AN222X1 g64168(.A (n_2159), .B (n_4778), .C (n_2160), .D (n_4774), .E
       (n_2164), .F (n_4779), .Q (n_6755));
  ON21X1 g64169(.A (n_3237), .B (n_1723), .C (n_5), .Q (n_6756));
  NA6I1X4 g64170(.B (n_3801), .C (n_3787), .D (n_4422), .E (n_6711), .F
       (n_6713), .AN (n_4202), .Q (n_6757));
  NO6I3X2 g64171(.D (n_4206), .E (n_3789), .F (n_3790), .AN (n_4203),
       .BN (n_3773), .CN (n_3774), .Q (n_6758));
  AN222X1 g64172(.A (n_3518), .B (n_4559), .C (n_3517), .D (n_4560), .E
       (n_3520), .F (n_4553), .Q (n_6759));
  AND4X2 g64173(.A (n_2426), .B (n_6786), .C (n_2424), .D (n_2425), .Q
       (n_6760));
  AN21X1 g64174(.A (n_272), .B (n_4466), .C (n_6761), .Q (n_6762));
  NA3X1 g64175(.A (n_679), .B (n_590), .C (n_649), .Q (n_6761));
  AN21X1 g64176(.A (n_272), .B (n_4461), .C (n_6763), .Q (n_6764));
  NA3X1 g64177(.A (n_656), .B (n_589), .C (n_627), .Q (n_6763));
  AN21X1 g64178(.A (n_272), .B (\rs1_data[26]_39276 ), .C (n_6765), .Q
       (n_6766));
  NA3X1 g64179(.A (n_670), .B (n_585), .C (n_635), .Q (n_6765));
  DFRQX1 \program_counter_reg[2] (.C (rc_gclk_205490), .D (n_434), .Q
       (program_counter[2]));
  DFRQX1 \program_counter_reg[3] (.C (rc_gclk_205490), .D (n_433), .Q
       (program_counter[3]));
  DFRQX1 \program_counter_reg[4] (.C (rc_gclk_205490), .D (n_435), .Q
       (program_counter[4]));
  DFRQX1 \program_counter_reg[5] (.C (rc_gclk_205490), .D (n_425), .Q
       (program_counter[5]));
  DFRQX1 \program_counter_reg[7] (.C (rc_gclk_205490), .D (n_437), .Q
       (program_counter[7]));
  DFRQX1 \program_counter_reg[6] (.C (rc_gclk_205490), .D (n_436), .Q
       (program_counter[6]));
  DFRQX1 \program_counter_reg[8] (.C (rc_gclk_205490), .D (n_430), .Q
       (program_counter[8]));
  DFRQX1 \program_counter_reg[9] (.C (rc_gclk_205490), .D (n_426), .Q
       (program_counter[9]));
  DFRQX1 \program_counter_reg[11] (.C (rc_gclk_205490), .D (n_427), .Q
       (program_counter[11]));
  DFRQX1 \program_counter_reg[10] (.C (rc_gclk_205490), .D (n_423), .Q
       (program_counter[10]));
  DFRQX1 \program_counter_reg[12] (.C (rc_gclk_205490), .D (n_418), .Q
       (program_counter[12]));
  DFRQX1 \program_counter_reg[13] (.C (rc_gclk_205490), .D (n_429), .Q
       (program_counter[13]));
  DFRQX1 \program_counter_reg[15] (.C (rc_gclk_205490), .D (n_422), .Q
       (program_counter[15]));
  DFRQX1 \program_counter_reg[14] (.C (rc_gclk_205490), .D (n_420), .Q
       (program_counter[14]));
  DFRQX1 \program_counter_reg[16] (.C (rc_gclk_205490), .D (n_421), .Q
       (program_counter[16]));
  DFRQX1 \program_counter_reg[17] (.C (rc_gclk_205490), .D (n_408), .Q
       (program_counter[17]));
  DFRQX1 \program_counter_reg[19] (.C (rc_gclk_205490), .D (n_416), .Q
       (program_counter[19]));
  DFRQX1 \program_counter_reg[18] (.C (rc_gclk_205490), .D (n_413), .Q
       (program_counter[18]));
  DFRQX1 \program_counter_reg[20] (.C (rc_gclk_205490), .D (n_414), .Q
       (program_counter[20]));
  DFRQX1 \program_counter_reg[21] (.C (rc_gclk_205490), .D (n_412), .Q
       (program_counter[21]));
  DFRQX1 \program_counter_reg[23] (.C (rc_gclk_205490), .D (n_415), .Q
       (program_counter[23]));
  DFRQX1 \program_counter_reg[22] (.C (rc_gclk_205490), .D (n_417), .Q
       (program_counter[22]));
  DFRQX1 \program_counter_reg[24] (.C (rc_gclk_205490), .D (n_407), .Q
       (program_counter[24]));
  DFRQX1 \program_counter_reg[25] (.C (rc_gclk_205490), .D (n_419), .Q
       (program_counter[25]));
  DFRQX1 \program_counter_reg[27] (.C (rc_gclk_205490), .D (n_431), .Q
       (program_counter[27]));
  DFRQX1 \program_counter_reg[26] (.C (rc_gclk_205490), .D (n_424), .Q
       (program_counter[26]));
  DFRQX1 \program_counter_reg[28] (.C (rc_gclk_205490), .D (n_428), .Q
       (program_counter[28]));
  DFRQX1 \program_counter_reg[29] (.C (rc_gclk_205490), .D (n_409), .Q
       (program_counter[29]));
  DFRQX1 \program_counter_reg[30] (.C (rc_gclk_205490), .D (n_410), .Q
       (program_counter[30]));
  DFRQX1 \program_counter_reg[31] (.C (rc_gclk_205490), .D (n_411), .Q
       (program_counter[31]));
  DFRQX1 \csr_mcause_code_reg[2] (.C (rc_gclk_205603), .D (n_10), .Q
       (csr_mcause_code[2]));
  DFRQX1 \csr_mcause_code_reg[4] (.C (rc_gclk_205603), .D (n_5627), .Q
       (csr_mcause_code[4]));
  DFRQX1 csr_mstatus_mie_reg(.C (rc_gclk), .D (n_940), .Q (n_5542));
  DFRQX1 \csr_mcycle_reg[32] (.C (clock), .D (n_1233), .Q
       (csr_mcycle[32]));
  DFRQX1 \csr_minstret_reg[32] (.C (rc_gclk), .D (n_1234), .Q
       (csr_minstret[32]));
  DFRQX1 \csr_mcycle_reg[42] (.C (clock), .D (n_1296), .Q
       (csr_mcycle[42]));
  DFRQX1 \csr_minstret_reg[42] (.C (rc_gclk), .D (n_1263), .Q
       (csr_minstret[42]));
  DFRQX1 \csr_mcycle_reg[44] (.C (clock), .D (n_1246), .Q
       (csr_mcycle[44]));
  DFRQX1 \csr_mcycle_reg[45] (.C (clock), .D (n_1255), .Q
       (csr_mcycle[45]));
  DFRQX1 \csr_mcycle_reg[46] (.C (clock), .D (n_1267), .Q
       (csr_mcycle[46]));
  DFRQX1 \csr_mcycle_reg[48] (.C (clock), .D (n_1245), .Q
       (csr_mcycle[48]));
  DFRQX1 \csr_minstret_reg[16] (.C (rc_gclk), .D (n_1195), .Q
       (csr_minstret[16]));
  DFRQX1 \csr_minstret_reg[17] (.C (rc_gclk), .D (n_1202), .Q
       (csr_minstret[17]));
  DFRQX1 \csr_mcycle_reg[49] (.C (clock), .D (n_1259), .Q
       (csr_mcycle[49]));
  DFRQX1 \csr_minstret_reg[50] (.C (rc_gclk), .D (n_1270), .Q
       (csr_minstret[50]));
  DFRQX1 \csr_mcycle_reg[50] (.C (clock), .D (n_1266), .Q
       (csr_mcycle[50]));
  DFRQX1 \csr_mcycle_reg[33] (.C (clock), .D (n_1236), .Q
       (csr_mcycle[33]));
  DFRQX1 \csr_minstret_reg[53] (.C (rc_gclk), .D (n_1269), .Q
       (csr_minstret[53]));
  DFRQX1 \csr_mcycle_reg[53] (.C (clock), .D (n_1265), .Q
       (csr_mcycle[53]));
  DFRQX1 \csr_mcycle_reg[54] (.C (clock), .D (n_1274), .Q
       (csr_mcycle[54]));
  DFRQX1 \csr_mcycle_reg[57] (.C (clock), .D (n_1278), .Q
       (csr_mcycle[57]));
  DFRQX1 \csr_mcycle_reg[61] (.C (clock), .D (n_1289), .Q
       (csr_mcycle[61]));
  DFRQX1 \csr_mcycle_reg[34] (.C (clock), .D (n_1241), .Q
       (csr_mcycle[34]));
  DFRQX1 \csr_mcycle_reg[36] (.C (clock), .D (n_1235), .Q
       (csr_mcycle[36]));
  DFRQX1 \csr_mcycle_reg[37] (.C (clock), .D (n_1240), .Q
       (csr_mcycle[37]));
  DFRQX1 \csr_mcycle_reg[38] (.C (clock), .D (n_1248), .Q
       (csr_mcycle[38]));
  DFRQX1 \csr_minstret_reg[38] (.C (rc_gclk), .D (n_1250), .Q
       (csr_minstret[38]));
  DFRQX1 \csr_mcycle_reg[40] (.C (clock), .D (n_1239), .Q
       (csr_mcycle[40]));
  DFRQX1 \csr_minstret_reg[40] (.C (rc_gclk), .D (n_1244), .Q
       (csr_minstret[40]));
  DFRQX1 \csr_mcycle_reg[41] (.C (clock), .D (n_1247), .Q
       (csr_mcycle[41]));
  DFRQX1 \csr_minstret_reg[41] (.C (rc_gclk), .D (n_1254), .Q
       (csr_minstret[41]));
  AND2X1 g64321(.A (n_2415), .B (n_2412), .Q (n_2799));
  AND2X1 g64323(.A (n_2438), .B (n_2442), .Q (n_2833));
  AND2X1 g64325(.A (n_3501), .B (n_3293), .Q (n_3516));
  AND6X1 g64327(.A (n_3823), .B (n_3824), .C (n_3831), .D (n_3832), .E
       (n_3316), .F (n_3311), .Q (n_6632));
  AND6X1 g64329(.A (n_6651), .B (n_4253), .C (n_3987), .D (n_4002), .E
       (n_3986), .F (n_4003), .Q (n_4451));
  AND2X2 g64331(.A (n_2078), .B (n_1949), .Q (n_2176));
  ON21X2 g64333(.A (n_2381), .B (n_3040), .C (n_3182), .Q
       (write_data[31]));
  ON21X2 g64335(.A (n_2381), .B (n_1643), .C (n_3181), .Q
       (write_data[30]));
  ON21X2 g64337(.A (n_2381), .B (n_3038), .C (n_3180), .Q
       (write_data[29]));
  ON21X2 g64339(.A (n_2381), .B (n_3042), .C (n_3179), .Q
       (write_data[28]));
  ON21X2 g64341(.A (n_2381), .B (n_3035), .C (n_3177), .Q
       (write_data[27]));
  ON21X2 g64343(.A (n_2381), .B (n_3044), .C (n_3183), .Q
       (write_data[26]));
  ON21X2 g64345(.A (n_2381), .B (n_6729), .C (n_3170), .Q
       (write_data[25]));
  ON21X2 g64347(.A (n_2381), .B (n_3032), .C (n_3178), .Q
       (write_data[24]));
  INX1 g64349(.A (take_trap_39145), .Q (n_175));
  INX2 g64351(.A (n_3483), .Q (n_3484));
  INX2 g64353(.A (n_1839), .Q (n_1838));
  INX2 g64355(.A (instruction[22]), .Q (n_1578));
  INX2 g64357(.A (n_1580), .Q (instruction[21]));
  INX2 g64359(.A (n_6787), .Q (n_1908));
  INX2 g64363(.A (n_3221), .Q (n_3220));
  AND2X4 g64364(.A (n_3500), .B (n_3487), .Q (n_6767));
  AND2X4 g64365(.A (n_3500), .B (n_3291), .Q (n_6768));
  AN221X1 g64373(.A (n_3295), .B (n_5184), .C (n_3505), .D (n_5170), .E
       (n_4192), .Q (n_6776));
  AN221X1 g64374(.A (n_3305), .B (n_4592), .C (n_3526), .D (n_4585), .E
       (n_4164), .Q (n_6777));
  AN221X1 g64375(.A (n_3296), .B (n_5091), .C (n_3505), .D (n_5077), .E
       (n_4099), .Q (n_6778));
  AN221X0 g64376(.A (n_3509), .B (n_5052), .C (n_3305), .D (n_5057), .E
       (n_4072), .Q (n_6779));
  AN221X1 g64377(.A (n_3538), .B (n_5284), .C (n_3540), .D (n_5285), .E
       (n_3900), .Q (n_6780));
  AN221X1 g64378(.A (n_3547), .B (n_5044), .C (n_3504), .D (n_5045), .E
       (n_3825), .Q (n_6781));
  AN222X0 g64379(.A (n_3520), .B (n_4925), .C (n_3518), .D (n_4931), .E
       (n_3517), .F (n_4932), .Q (n_6782));
  AN21X1 g64380(.A (n_3520), .B (n_4677), .C (n_3879), .Q (n_6783));
  AN222X0 g64381(.A (n_3518), .B (n_5024), .C (n_3517), .D (n_5025), .E
       (n_3520), .F (n_5018), .Q (n_6784));
  ON221X1 g64382(.A (n_1594), .B (n_1707), .C (n_2189), .D (n_1705), .E
       (n_2541), .Q (n_6785));
  AN21X1 g64383(.A (n_1813), .B (n_4890), .C (n_2294), .Q (n_6786));
  AO21X4 g64384(.A (n_1725), .B (instruction[22]), .C (n_1764), .Q
       (n_6787));
  DFRQX1 \csr_mcause_code_reg[3] (.C (rc_gclk_205603), .D (n_9), .Q
       (csr_mcause_code[3]));
  DFRQX1 \csr_mcause_code_reg[1] (.C (rc_gclk_205603), .D (n_12), .Q
       (csr_mcause_code[1]));
  DFRQX1 \csr_mcause_code_reg[0] (.C (rc_gclk_205603), .D (n_14), .Q
       (csr_mcause_code[0]));
  DFRQX1 \csr_minstret_reg[20] (.C (rc_gclk), .D (n_1201), .Q
       (csr_minstret[20]));
  DFRQX1 \csr_mcycle_reg[52] (.C (clock), .D (n_1258), .Q
       (csr_mcycle[52]));
  AND2X1 g64396(.A (n_2411), .B (n_2405), .Q (n_2808));
  AND6X1 g64400(.A (n_1621), .B (n_2848), .C (n_2856), .D (n_2855), .E
       (n_2585), .F (n_2475), .Q (n_3038));
  INX2 g64402(.A (\instruction[14]_40077 ), .Q (n_1687));
  INX1 g64404(.A (n_1661), .Q (take_trap_39145));
endmodule

