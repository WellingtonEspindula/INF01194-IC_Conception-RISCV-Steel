
module iopads(clock, reset, halt, 
	rw_address,
	read_data,
	read_request,
	read_response,
	write_data,
	write_strobe,
	write_request,
	write_response,
	irq_external,
	irq_external_response,
	irq_timer,
	irq_timer_response,
	irq_software,
	irq_software_response,
	irq_fast,
	irq_fast_response,
	real_time_clock,
     rw_address_O,
     clock_I, reset_I, halt_I,
     read_data_I,
     read_request_O,
     read_response_I,
     write_data_O,
     write_strobe_O,
     write_request_O,
     write_response_I,
     irq_external_I,
     irq_external_response_O,
     irq_timer_I,
     irq_timer_response_O,
     irq_software_I,
     irq_software_response_O,
     irq_fast_I,
     irq_fast_response_O,
     real_time_clock_I);

     input clock, reset, halt;
	output [31:0] rw_address;
	input [31:0] read_data;
	output read_request;
	input read_response;
	output [31:0] write_data;
	output [3:0] write_strobe;
	output write_request;
     input write_response;
     input irq_external;
	output irq_external_response;
	input irq_timer;
	output irq_timer_response;
	input irq_software;
	output irq_software_response;
	input [15:0] irq_fast;
	output [15:0] irq_fast_response;
     input  [63:0] real_time_clock;

     output clock_I, reset_I, halt_I;
     input [31:0]  rw_address_O;
     output  [31:0]  read_data_I;
     input read_request_O;
     output  read_response_I;
     input [31:0]  write_data_O;
     input [3:0 ]  write_strobe_O;
     input write_request_O;
     output  write_response_I;
     output  irq_external_I;
     input irq_external_response_O;
     output  irq_timer_I;
     input irq_timer_response_O;
     output  irq_software_I;
     input irq_software_response_O;
     output  [15:0]  irq_fast_I;
     input [15:0]  irq_fast_response_O;
     output  [63:0]  real_time_clock_I;

     ICP PAD_clk_i(.PAD(clock), .Y(clock_I));
     ICP PAD_reset_i(.PAD(reset), .Y(reset_I));
     ICP PAD_halt_i(.PAD(halt), .Y(halt_I));

     BD8P PAD_rw_address_o_0(.A(rw_address_O[0]), .PAD(rw_address[0]));
     BD8P PAD_rw_address_o_1(.A(rw_address_O[1]), .PAD(rw_address[1]));
     BD8P PAD_rw_address_o_2(.A(rw_address_O[2]), .PAD(rw_address[2]));
     BD8P PAD_rw_address_o_3(.A(rw_address_O[3]), .PAD(rw_address[3]));
     BD8P PAD_rw_address_o_4(.A(rw_address_O[4]), .PAD(rw_address[4]));
     BD8P PAD_rw_address_o_5(.A(rw_address_O[5]), .PAD(rw_address[5]));
     BD8P PAD_rw_address_o_6(.A(rw_address_O[6]), .PAD(rw_address[6]));
     BD8P PAD_rw_address_o_7(.A(rw_address_O[7]), .PAD(rw_address[7]));
     BD8P PAD_rw_address_o_8(.A(rw_address_O[8]), .PAD(rw_address[8]));
     BD8P PAD_rw_address_o_9(.A(rw_address_O[9]), .PAD(rw_address[9]));
     BD8P PAD_rw_address_o_10(.A(rw_address_O[10]), .PAD(rw_address[10]));
     BD8P PAD_rw_address_o_11(.A(rw_address_O[11]), .PAD(rw_address[11]));
     BD8P PAD_rw_address_o_12(.A(rw_address_O[12]), .PAD(rw_address[12]));
     BD8P PAD_rw_address_o_13(.A(rw_address_O[13]), .PAD(rw_address[13]));
     BD8P PAD_rw_address_o_14(.A(rw_address_O[14]), .PAD(rw_address[14]));
     BD8P PAD_rw_address_o_15(.A(rw_address_O[15]), .PAD(rw_address[15]));
     BD8P PAD_rw_address_o_16(.A(rw_address_O[16]), .PAD(rw_address[16]));
     BD8P PAD_rw_address_o_17(.A(rw_address_O[17]), .PAD(rw_address[17]));
     BD8P PAD_rw_address_o_18(.A(rw_address_O[18]), .PAD(rw_address[18]));
     BD8P PAD_rw_address_o_19(.A(rw_address_O[19]), .PAD(rw_address[19]));
     BD8P PAD_rw_address_o_20(.A(rw_address_O[20]), .PAD(rw_address[20]));
     BD8P PAD_rw_address_o_21(.A(rw_address_O[21]), .PAD(rw_address[21]));
     BD8P PAD_rw_address_o_22(.A(rw_address_O[22]), .PAD(rw_address[22]));
     BD8P PAD_rw_address_o_23(.A(rw_address_O[23]), .PAD(rw_address[23]));
     BD8P PAD_rw_address_o_24(.A(rw_address_O[24]), .PAD(rw_address[24]));
     BD8P PAD_rw_address_o_25(.A(rw_address_O[25]), .PAD(rw_address[25]));
     BD8P PAD_rw_address_o_26(.A(rw_address_O[26]), .PAD(rw_address[26]));
     BD8P PAD_rw_address_o_27(.A(rw_address_O[27]), .PAD(rw_address[27]));
     BD8P PAD_rw_address_o_28(.A(rw_address_O[28]), .PAD(rw_address[28]));
     BD8P PAD_rw_address_o_29(.A(rw_address_O[29]), .PAD(rw_address[29]));
     BD8P PAD_rw_address_o_30(.A(rw_address_O[30]), .PAD(rw_address[30]));
     BD8P PAD_rw_address_o_31(.A(rw_address_O[31]), .PAD(rw_address[31]));

     ICP PAD_read_data_i_0(.PAD(read_data[0]), .Y(read_data_I[0]));
     ICP PAD_read_data_i_1(.PAD(read_data[1]), .Y(read_data_I[1]));
     ICP PAD_read_data_i_2(.PAD(read_data[2]), .Y(read_data_I[2]));
     ICP PAD_read_data_i_3(.PAD(read_data[3]), .Y(read_data_I[3]));
     ICP PAD_read_data_i_4(.PAD(read_data[4]), .Y(read_data_I[4]));
     ICP PAD_read_data_i_5(.PAD(read_data[5]), .Y(read_data_I[5]));
     ICP PAD_read_data_i_6(.PAD(read_data[6]), .Y(read_data_I[6]));
     ICP PAD_read_data_i_7(.PAD(read_data[7]), .Y(read_data_I[7]));
     ICP PAD_read_data_i_8(.PAD(read_data[8]), .Y(read_data_I[8]));
     ICP PAD_read_data_i_9(.PAD(read_data[9]), .Y(read_data_I[9]));
     ICP PAD_read_data_i_10(.PAD(read_data[10]), .Y(read_data_I[10]));
     ICP PAD_read_data_i_11(.PAD(read_data[11]), .Y(read_data_I[11]));
     ICP PAD_read_data_i_12(.PAD(read_data[12]), .Y(read_data_I[12]));
     ICP PAD_read_data_i_13(.PAD(read_data[13]), .Y(read_data_I[13]));
     ICP PAD_read_data_i_14(.PAD(read_data[14]), .Y(read_data_I[14]));
     ICP PAD_read_data_i_15(.PAD(read_data[15]), .Y(read_data_I[15]));
     ICP PAD_read_data_i_16(.PAD(read_data[16]), .Y(read_data_I[16]));
     ICP PAD_read_data_i_17(.PAD(read_data[17]), .Y(read_data_I[17]));
     ICP PAD_read_data_i_18(.PAD(read_data[18]), .Y(read_data_I[18]));
     ICP PAD_read_data_i_19(.PAD(read_data[19]), .Y(read_data_I[19]));
     ICP PAD_read_data_i_20(.PAD(read_data[20]), .Y(read_data_I[20]));
     ICP PAD_read_data_i_21(.PAD(read_data[21]), .Y(read_data_I[21]));
     ICP PAD_read_data_i_22(.PAD(read_data[22]), .Y(read_data_I[22]));
     ICP PAD_read_data_i_23(.PAD(read_data[23]), .Y(read_data_I[23]));
     ICP PAD_read_data_i_24(.PAD(read_data[24]), .Y(read_data_I[24]));
     ICP PAD_read_data_i_25(.PAD(read_data[25]), .Y(read_data_I[25]));
     ICP PAD_read_data_i_26(.PAD(read_data[26]), .Y(read_data_I[26]));
     ICP PAD_read_data_i_27(.PAD(read_data[27]), .Y(read_data_I[27]));
     ICP PAD_read_data_i_28(.PAD(read_data[28]), .Y(read_data_I[28]));
     ICP PAD_read_data_i_29(.PAD(read_data[29]), .Y(read_data_I[29]));
     ICP PAD_read_data_i_30(.PAD(read_data[30]), .Y(read_data_I[30]));
     ICP PAD_read_data_i_31(.PAD(read_data[31]), .Y(read_data_I[31]));

     BD8P PAD_read_request_o(.A(read_request_O), .PAD(read_request));
     ICP PAD_read_response_i(.PAD(read_response), .Y(read_response_I));

     BD8P PAD_write_data_o_0(.A(write_data_O[0]), .PAD(write_data[0]));
     BD8P PAD_write_data_o_1(.A(write_data_O[1]), .PAD(write_data[1]));
     BD8P PAD_write_data_o_2(.A(write_data_O[2]), .PAD(write_data[2]));
     BD8P PAD_write_data_o_3(.A(write_data_O[3]), .PAD(write_data[3]));
     BD8P PAD_write_data_o_4(.A(write_data_O[4]), .PAD(write_data[4]));
     BD8P PAD_write_data_o_5(.A(write_data_O[5]), .PAD(write_data[5]));
     BD8P PAD_write_data_o_6(.A(write_data_O[6]), .PAD(write_data[6]));
     BD8P PAD_write_data_o_7(.A(write_data_O[7]), .PAD(write_data[7]));
     BD8P PAD_write_data_o_8(.A(write_data_O[8]), .PAD(write_data[8]));
     BD8P PAD_write_data_o_9(.A(write_data_O[9]), .PAD(write_data[9]));
     BD8P PAD_write_data_o_10(.A(write_data_O[10]), .PAD(write_data[10]));
     BD8P PAD_write_data_o_11(.A(write_data_O[11]), .PAD(write_data[11]));
     BD8P PAD_write_data_o_12(.A(write_data_O[12]), .PAD(write_data[12]));
     BD8P PAD_write_data_o_13(.A(write_data_O[13]), .PAD(write_data[13]));
     BD8P PAD_write_data_o_14(.A(write_data_O[14]), .PAD(write_data[14]));
     BD8P PAD_write_data_o_15(.A(write_data_O[15]), .PAD(write_data[15]));
     BD8P PAD_write_data_o_16(.A(write_data_O[16]), .PAD(write_data[16]));
     BD8P PAD_write_data_o_17(.A(write_data_O[17]), .PAD(write_data[17]));
     BD8P PAD_write_data_o_18(.A(write_data_O[18]), .PAD(write_data[18]));
     BD8P PAD_write_data_o_19(.A(write_data_O[19]), .PAD(write_data[19]));
     BD8P PAD_write_data_o_20(.A(write_data_O[20]), .PAD(write_data[20]));
     BD8P PAD_write_data_o_21(.A(write_data_O[21]), .PAD(write_data[21]));
     BD8P PAD_write_data_o_22(.A(write_data_O[22]), .PAD(write_data[22]));
     BD8P PAD_write_data_o_23(.A(write_data_O[23]), .PAD(write_data[23]));
     BD8P PAD_write_data_o_24(.A(write_data_O[24]), .PAD(write_data[24]));
     BD8P PAD_write_data_o_25(.A(write_data_O[25]), .PAD(write_data[25]));
     BD8P PAD_write_data_o_26(.A(write_data_O[26]), .PAD(write_data[26]));
     BD8P PAD_write_data_o_27(.A(write_data_O[27]), .PAD(write_data[27]));
     BD8P PAD_write_data_o_28(.A(write_data_O[28]), .PAD(write_data[28]));
     BD8P PAD_write_data_o_29(.A(write_data_O[29]), .PAD(write_data[29]));
     BD8P PAD_write_data_o_30(.A(write_data_O[30]), .PAD(write_data[30]));
     BD8P PAD_write_data_o_31(.A(write_data_O[31]), .PAD(write_data[31]));

     BD8P PAD_write_strobe_o_0(.A(write_strobe_O[0]), .PAD(write_strobe[0]));
     BD8P PAD_write_strobe_o_1(.A(write_strobe_O[1]), .PAD(write_strobe[1]));
     BD8P PAD_write_strobe_o_2(.A(write_strobe_O[2]), .PAD(write_strobe[2]));
     BD8P PAD_write_strobe_o_3(.A(write_strobe_O[3]), .PAD(write_strobe[3]));
     
     BD8P PAD_write_request_o(.A(write_request_O), .PAD(write_request));
     ICP PAD_write_response_i(.PAD(write_response), .Y(write_response_I));

     ICP PAD_irq_external_i(.PAD(irq_external), .Y(irq_external_I));
     BD8P PAD_irq_external_response_o(.A(irq_external_response_O), .PAD(irq_external_response));

     ICP PAD_irq_timer_i(.PAD(irq_timer), .Y(irq_timer_I));
     BD8P PAD_irq_timer_response_o(.A(irq_timer_response_O), .PAD(irq_timer_response));

     ICP PAD_irq_software_i(.PAD(irq_software), .Y(irq_software_I));
     BD8P PAD_irq_software_response_o(.A(irq_software_response_O), .PAD(irq_software_response));
     
     ICP PAD_irq_fast_i_0(.PAD(irq_fast[0]), .Y(irq_fast_I[0]));
     ICP PAD_irq_fast_i_1(.PAD(irq_fast[1]), .Y(irq_fast_I[1]));
     ICP PAD_irq_fast_i_2(.PAD(irq_fast[2]), .Y(irq_fast_I[2]));
     ICP PAD_irq_fast_i_3(.PAD(irq_fast[3]), .Y(irq_fast_I[3]));
     ICP PAD_irq_fast_i_4(.PAD(irq_fast[4]), .Y(irq_fast_I[4]));
     ICP PAD_irq_fast_i_5(.PAD(irq_fast[5]), .Y(irq_fast_I[5]));
     ICP PAD_irq_fast_i_6(.PAD(irq_fast[6]), .Y(irq_fast_I[6]));
     ICP PAD_irq_fast_i_7(.PAD(irq_fast[7]), .Y(irq_fast_I[7]));
     ICP PAD_irq_fast_i_8(.PAD(irq_fast[8]), .Y(irq_fast_I[8]));
     ICP PAD_irq_fast_i_9(.PAD(irq_fast[9]), .Y(irq_fast_I[9]));
     ICP PAD_irq_fast_i_10(.PAD(irq_fast[10]), .Y(irq_fast_I[10]));
     ICP PAD_irq_fast_i_11(.PAD(irq_fast[11]), .Y(irq_fast_I[11]));
     ICP PAD_irq_fast_i_12(.PAD(irq_fast[12]), .Y(irq_fast_I[12]));
     ICP PAD_irq_fast_i_13(.PAD(irq_fast[13]), .Y(irq_fast_I[13]));
     ICP PAD_irq_fast_i_14(.PAD(irq_fast[14]), .Y(irq_fast_I[14]));
     ICP PAD_irq_fast_i_15(.PAD(irq_fast[15]), .Y(irq_fast_I[15]));

     BD8P PAD_irq_fast_response_o_0(.A(irq_fast_response_O[0]), .PAD(irq_fast_response[0]));
     BD8P PAD_irq_fast_response_o_1(.A(irq_fast_response_O[1]), .PAD(irq_fast_response[1]));
     BD8P PAD_irq_fast_response_o_2(.A(irq_fast_response_O[2]), .PAD(irq_fast_response[2]));
     BD8P PAD_irq_fast_response_o_3(.A(irq_fast_response_O[3]), .PAD(irq_fast_response[3]));
     BD8P PAD_irq_fast_response_o_4(.A(irq_fast_response_O[4]), .PAD(irq_fast_response[4]));
     BD8P PAD_irq_fast_response_o_5(.A(irq_fast_response_O[5]), .PAD(irq_fast_response[5]));
     BD8P PAD_irq_fast_response_o_6(.A(irq_fast_response_O[6]), .PAD(irq_fast_response[6]));
     BD8P PAD_irq_fast_response_o_7(.A(irq_fast_response_O[7]), .PAD(irq_fast_response[7]));
     BD8P PAD_irq_fast_response_o_8(.A(irq_fast_response_O[8]), .PAD(irq_fast_response[8]));
     BD8P PAD_irq_fast_response_o_9(.A(irq_fast_response_O[9]), .PAD(irq_fast_response[9]));
     BD8P PAD_irq_fast_response_o_10(.A(irq_fast_response_O[10]), .PAD(irq_fast_response[10]));
     BD8P PAD_irq_fast_response_o_11(.A(irq_fast_response_O[11]), .PAD(irq_fast_response[11]));
     BD8P PAD_irq_fast_response_o_12(.A(irq_fast_response_O[12]), .PAD(irq_fast_response[12]));
     BD8P PAD_irq_fast_response_o_13(.A(irq_fast_response_O[13]), .PAD(irq_fast_response[13]));
     BD8P PAD_irq_fast_response_o_14(.A(irq_fast_response_O[14]), .PAD(irq_fast_response[14]));
     BD8P PAD_irq_fast_response_o_15(.A(irq_fast_response_O[15]), .PAD(irq_fast_response[15]));

     ICP PAD_real_time_clock_i_0(.PAD(real_time_clock[0]), .Y(real_time_clock_I[0]));
     ICP PAD_real_time_clock_i_1(.PAD(real_time_clock[1]), .Y(real_time_clock_I[1]));
     ICP PAD_real_time_clock_i_2(.PAD(real_time_clock[2]), .Y(real_time_clock_I[2]));
     ICP PAD_real_time_clock_i_3(.PAD(real_time_clock[3]), .Y(real_time_clock_I[3]));
     ICP PAD_real_time_clock_i_4(.PAD(real_time_clock[4]), .Y(real_time_clock_I[4]));
     ICP PAD_real_time_clock_i_5(.PAD(real_time_clock[5]), .Y(real_time_clock_I[5]));
     ICP PAD_real_time_clock_i_6(.PAD(real_time_clock[6]), .Y(real_time_clock_I[6]));
     ICP PAD_real_time_clock_i_7(.PAD(real_time_clock[7]), .Y(real_time_clock_I[7]));
     ICP PAD_real_time_clock_i_8(.PAD(real_time_clock[8]), .Y(real_time_clock_I[8]));
     ICP PAD_real_time_clock_i_9(.PAD(real_time_clock[9]), .Y(real_time_clock_I[9]));
     ICP PAD_real_time_clock_i_10(.PAD(real_time_clock[10]), .Y(real_time_clock_I[10]));
     ICP PAD_real_time_clock_i_11(.PAD(real_time_clock[11]), .Y(real_time_clock_I[11]));
     ICP PAD_real_time_clock_i_12(.PAD(real_time_clock[12]), .Y(real_time_clock_I[12]));
     ICP PAD_real_time_clock_i_13(.PAD(real_time_clock[13]), .Y(real_time_clock_I[13]));
     ICP PAD_real_time_clock_i_14(.PAD(real_time_clock[14]), .Y(real_time_clock_I[14]));
     ICP PAD_real_time_clock_i_15(.PAD(real_time_clock[15]), .Y(real_time_clock_I[15]));
     ICP PAD_real_time_clock_i_16(.PAD(real_time_clock[16]), .Y(real_time_clock_I[16]));
     ICP PAD_real_time_clock_i_17(.PAD(real_time_clock[17]), .Y(real_time_clock_I[17]));
     ICP PAD_real_time_clock_i_18(.PAD(real_time_clock[18]), .Y(real_time_clock_I[18]));
     ICP PAD_real_time_clock_i_19(.PAD(real_time_clock[19]), .Y(real_time_clock_I[19]));
     ICP PAD_real_time_clock_i_20(.PAD(real_time_clock[20]), .Y(real_time_clock_I[20]));
     ICP PAD_real_time_clock_i_21(.PAD(real_time_clock[21]), .Y(real_time_clock_I[21]));
     ICP PAD_real_time_clock_i_22(.PAD(real_time_clock[22]), .Y(real_time_clock_I[22]));
     ICP PAD_real_time_clock_i_23(.PAD(real_time_clock[23]), .Y(real_time_clock_I[23]));
     ICP PAD_real_time_clock_i_24(.PAD(real_time_clock[24]), .Y(real_time_clock_I[24]));
     ICP PAD_real_time_clock_i_25(.PAD(real_time_clock[25]), .Y(real_time_clock_I[25]));
     ICP PAD_real_time_clock_i_26(.PAD(real_time_clock[26]), .Y(real_time_clock_I[26]));
     ICP PAD_real_time_clock_i_27(.PAD(real_time_clock[27]), .Y(real_time_clock_I[27]));
     ICP PAD_real_time_clock_i_28(.PAD(real_time_clock[28]), .Y(real_time_clock_I[28]));
     ICP PAD_real_time_clock_i_29(.PAD(real_time_clock[29]), .Y(real_time_clock_I[29]));
     ICP PAD_real_time_clock_i_30(.PAD(real_time_clock[30]), .Y(real_time_clock_I[30]));
     ICP PAD_real_time_clock_i_31(.PAD(real_time_clock[31]), .Y(real_time_clock_I[31]));
     ICP PAD_real_time_clock_i_32(.PAD(real_time_clock[32]), .Y(real_time_clock_I[32]));
     ICP PAD_real_time_clock_i_33(.PAD(real_time_clock[33]), .Y(real_time_clock_I[33]));
     ICP PAD_real_time_clock_i_34(.PAD(real_time_clock[34]), .Y(real_time_clock_I[34]));
     ICP PAD_real_time_clock_i_35(.PAD(real_time_clock[35]), .Y(real_time_clock_I[35]));
     ICP PAD_real_time_clock_i_36(.PAD(real_time_clock[36]), .Y(real_time_clock_I[36]));
     ICP PAD_real_time_clock_i_37(.PAD(real_time_clock[37]), .Y(real_time_clock_I[37]));
     ICP PAD_real_time_clock_i_38(.PAD(real_time_clock[38]), .Y(real_time_clock_I[38]));
     ICP PAD_real_time_clock_i_39(.PAD(real_time_clock[39]), .Y(real_time_clock_I[39]));
     ICP PAD_real_time_clock_i_40(.PAD(real_time_clock[40]), .Y(real_time_clock_I[40]));
     ICP PAD_real_time_clock_i_41(.PAD(real_time_clock[41]), .Y(real_time_clock_I[41]));
     ICP PAD_real_time_clock_i_42(.PAD(real_time_clock[42]), .Y(real_time_clock_I[42]));
     ICP PAD_real_time_clock_i_43(.PAD(real_time_clock[43]), .Y(real_time_clock_I[43]));
     ICP PAD_real_time_clock_i_44(.PAD(real_time_clock[44]), .Y(real_time_clock_I[44]));
     ICP PAD_real_time_clock_i_45(.PAD(real_time_clock[45]), .Y(real_time_clock_I[45]));
     ICP PAD_real_time_clock_i_46(.PAD(real_time_clock[46]), .Y(real_time_clock_I[46]));
     ICP PAD_real_time_clock_i_47(.PAD(real_time_clock[47]), .Y(real_time_clock_I[47]));
     ICP PAD_real_time_clock_i_48(.PAD(real_time_clock[48]), .Y(real_time_clock_I[48]));
     ICP PAD_real_time_clock_i_49(.PAD(real_time_clock[49]), .Y(real_time_clock_I[49]));
     ICP PAD_real_time_clock_i_50(.PAD(real_time_clock[50]), .Y(real_time_clock_I[50]));
     ICP PAD_real_time_clock_i_51(.PAD(real_time_clock[51]), .Y(real_time_clock_I[51]));
     ICP PAD_real_time_clock_i_52(.PAD(real_time_clock[52]), .Y(real_time_clock_I[52]));
     ICP PAD_real_time_clock_i_53(.PAD(real_time_clock[53]), .Y(real_time_clock_I[53]));
     ICP PAD_real_time_clock_i_54(.PAD(real_time_clock[54]), .Y(real_time_clock_I[54]));
     ICP PAD_real_time_clock_i_55(.PAD(real_time_clock[55]), .Y(real_time_clock_I[55]));
     ICP PAD_real_time_clock_i_56(.PAD(real_time_clock[56]), .Y(real_time_clock_I[56]));
     ICP PAD_real_time_clock_i_57(.PAD(real_time_clock[57]), .Y(real_time_clock_I[57]));
     ICP PAD_real_time_clock_i_58(.PAD(real_time_clock[58]), .Y(real_time_clock_I[58]));
     ICP PAD_real_time_clock_i_59(.PAD(real_time_clock[59]), .Y(real_time_clock_I[59]));
     ICP PAD_real_time_clock_i_60(.PAD(real_time_clock[60]), .Y(real_time_clock_I[60]));
     ICP PAD_real_time_clock_i_61(.PAD(real_time_clock[61]), .Y(real_time_clock_I[61]));
     ICP PAD_real_time_clock_i_62(.PAD(real_time_clock[62]), .Y(real_time_clock_I[62]));
     ICP PAD_real_time_clock_i_63(.PAD(real_time_clock[63]), .Y(real_time_clock_I[63]));

	VDDORPADP PAD_vdd_E();
	VDDPADP PAD_vdd_core_E();

	VDDPADP PAD_vdd_core_N();
	GNDORPADP PAD_vss_core_N();

	GNDORPADP PAD_vss_W();

	GNDORPADP PAD_vss_S();

	CORNERP PAD_corner_ll();
	CORNERP PAD_corner_lr();
	CORNERP PAD_corner_ul();
	CORNERP PAD_corner_ur();	
endmodule

module top(clock, 
              reset, 
              halt, 
              rw_address,
              read_data,
              read_request,
              read_response,
              write_data,
              write_strobe,
              write_request,
              write_response,
              irq_external,
              irq_external_response,
              irq_timer,
              irq_timer_response,
              irq_software,
              irq_software_response,
              irq_fast,
              irq_fast_response,
              real_time_clock);

     input  clock;
     input  reset;
     input  halt;

     output [31:0]  rw_address;
     input [31:0]  read_data;
     output  read_request;
     input  read_response;
     output [31:0]  write_data;
     output [3:0 ]  write_strobe;
     output  write_request;
     input  write_response;

     input  irq_external;
     output  irq_external_response;
     input  irq_timer;
     output  irq_timer_response;
     input  irq_software;
     output  irq_software_response;
     input [15:0]  irq_fast;
     output [15:0]  irq_fast_response;

     input [63:0]  real_time_clock;


	wire clock_I, reset_I, halt_I;
	
	wire [31:0]  rw_address_O;
	wire  [31:0]  read_data_I;
	wire read_request_O;
	wire  read_response_I;
	wire [31:0]  write_data_O;
	wire [3:0 ]  write_strobe_O;
	wire write_request_O;

	wire  write_response_I;

	wire  irq_external_I;
	wire irq_external_response_O;
	wire  irq_timer_I;
	wire irq_timer_response_O;
	wire  irq_software_I;
	wire irq_software_response_O;
	wire  [15:0]  irq_fast_I;
	wire [15:0]  irq_fast_response_O;

	wire  [63:0]  real_time_clock_I;

	rvsteel_core top_INST(
		.clock(clock_I),
		.reset(reset_I),
          .halt(halt_I),
          .rw_address(rw_address_O),
          .read_data(read_data_I),
          .read_request(read_request_O),
          .read_response(read_response_I),
          .write_data(write_data_O),
          .write_strobe(write_strobe_O),
          .write_request(write_request_O),
          .write_response(write_response_I),
          .irq_external(irq_external_I),
          .irq_external_response(irq_external_response_O),
          .irq_timer(irq_timer_I),
          .irq_timer_response(irq_timer_response_O),
          .irq_software(irq_software_I),
          .irq_software_response(irq_software_response_O),
          .irq_fast(irq_fast_I),
          .irq_fast_response(irq_fast_response_O),
          .real_time_clock(real_time_clock_I)
	);

	iopads IOPADS_INST(
          .clock(clock),
          .reset(reset),
          .halt(halt),
          .rw_address(rw_address),
          .read_data(read_data),
          .read_request(read_request),
          .read_response(read_response),
          .write_data(write_data),
          .write_strobe(write_strobe),
          .write_request(write_request),
          .write_response(write_response),
          .irq_external(irq_external),
          .irq_external_response(irq_external_response),
          .irq_timer(irq_timer),
          .irq_timer_response(irq_timer_response),
          .irq_software(irq_software),
          .irq_software_response(irq_software_response),
          .irq_fast(irq_fast),
          .irq_fast_response(irq_fast_response),
          .real_time_clock(real_time_clock)
	);
endmodule



// Generated by Cadence Genus(TM) Synthesis Solution GENUS15.22 - 15.20-s024_1
// Generated on: Nov 13 2024 23:22:17

// Verification Directory fv/rvsteel_core 

module RC_CG_MOD_AUTO_rvsteel_core(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_9(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_10(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_11(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_12(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_13(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_14(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_15(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_16(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_17(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_18(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_1(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_19(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_20(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_21(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_22(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_23(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_7;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_7), .Q (enl));
  OR2X1 g13(.A (enable), .B (test), .Q (n_7));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_24(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_25(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_26(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_27(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_28(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_2(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_29(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_30(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_31(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_32(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_33(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_34(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_35(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_36(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_37(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_38(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_3(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_7;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_7), .Q (enl));
  OR2X1 g13(.A (enable), .B (test), .Q (n_7));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_39(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_7;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_7), .Q (enl));
  OR2X1 g13(.A (enable), .B (test), .Q (n_7));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_40(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_41(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_4(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_5(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_6(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_7(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module RC_CG_MOD_AUTO_rvsteel_core_8(ck_in, enable, test, ck_out);
  input ck_in, enable, test;
  output ck_out;
  wire ck_in, enable, test;
  wire ck_out;
  wire enl, n_0;
  AND2X1 g12(.A (ck_in), .B (enl), .Q (ck_out));
  DLLQX1 enl_reg(.GN (ck_in), .D (n_0), .Q (enl));
  OR2X1 g7(.A (enable), .B (test), .Q (n_0));
endmodule

module csa_tree_add_1660_20_group_293(in_0, in_1, in_2, out_0);
  input [31:0] in_0;
  input [33:0] in_1, in_2;
  output [31:0] out_0;
  wire [31:0] in_0;
  wire [33:0] in_1, in_2;
  wire [31:0] out_0;
  wire n_95, n_96, n_97, n_99, n_101, n_102, n_106, n_108;
  wire n_109, n_110, n_113, n_114, n_115, n_118, n_119, n_120;
  wire n_121, n_124, n_128, n_129, n_131, n_133, n_134, n_135;
  wire n_139, n_142, n_143, n_144, n_146, n_147, n_148, n_151;
  wire n_153, n_154, n_155, n_157, n_166, n_167, n_168, n_169;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_268, n_269, n_270, n_271;
  wire n_274, n_275, n_276, n_277, n_278, n_280, n_282, n_284;
  wire n_286, n_287, n_288, n_290, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_324;
  wire n_326, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_340, n_341, n_344, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
  wire n_382, n_383, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_432, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_464;
  HAX2 g251(.A (in_1[14]), .B (in_0[14]), .S (n_108), .CO (n_142));
  HAX2 g252(.A (in_1[24]), .B (in_0[24]), .S (n_119), .CO (n_153));
  HAX2 g253(.A (in_1[25]), .B (in_0[25]), .S (n_120), .CO (n_154));
  HAX2 g254(.A (in_1[26]), .B (in_0[26]), .S (n_121), .CO (n_155));
  HAX2 g258(.A (in_1[28]), .B (in_0[28]), .S (n_124), .CO (n_157));
  HAX2 g263(.A (in_1[2]), .B (in_0[2]), .S (n_95), .CO (n_128));
  HAX2 g264(.A (in_1[3]), .B (in_0[3]), .S (n_96), .CO (n_129));
  HAX2 g265(.A (in_1[15]), .B (in_0[15]), .S (n_109), .CO (n_143));
  HAX2 g266(.A (in_1[4]), .B (in_0[4]), .S (n_97), .CO (n_131));
  HAX2 g270(.A (in_1[6]), .B (in_0[6]), .S (n_99), .CO (n_133));
  HAX2 g271(.A (in_1[7]), .B (in_0[7]), .S (n_101), .CO (n_134));
  HAX2 g272(.A (in_1[8]), .B (in_0[8]), .S (n_102), .CO (n_135));
  HAX2 g282(.A (in_1[12]), .B (in_0[12]), .S (n_106), .CO (n_139));
  HAX2 g286(.A (in_1[16]), .B (in_0[16]), .S (n_110), .CO (n_144));
  HAX2 g290(.A (in_1[18]), .B (in_0[18]), .S (n_113), .CO (n_146));
  HAX2 g291(.A (in_1[19]), .B (in_0[19]), .S (n_114), .CO (n_147));
  HAX2 g292(.A (in_1[20]), .B (in_0[20]), .S (n_115), .CO (n_148));
  HAX2 g299(.A (in_1[23]), .B (in_0[23]), .S (n_118), .CO (n_151));
  EO2X1 g982(.A (n_399), .B (n_250), .Q (out_0[20]));
  EO2X1 g985(.A (n_411), .B (n_251), .Q (out_0[24]));
  EO2X1 g986(.A (n_410), .B (n_252), .Q (out_0[18]));
  EO2X1 g987(.A (n_409), .B (n_241), .Q (out_0[17]));
  AND2X4 g989(.A (n_401), .B (n_362), .Q (n_412));
  MU2IX1 g990(.S (n_246), .IN0 (n_395), .IN1 (n_394), .Q (out_0[16]));
  AN21X1 g991(.A (n_394), .B (n_330), .C (n_363), .Q (n_411));
  AN21X1 g992(.A (n_394), .B (n_257), .C (n_301), .Q (n_410));
  AN21X1 g993(.A (n_394), .B (n_179), .C (n_181), .Q (n_409));
  AN21X1 g994(.A (n_394), .B (n_347), .C (n_374), .Q (n_408));
  AN21X1 g995(.A (n_394), .B (n_351), .C (n_378), .Q (n_407));
  AN21X1 g996(.A (n_394), .B (n_354), .C (n_377), .Q (n_406));
  AN21X1 g997(.A (n_394), .B (n_328), .C (n_361), .Q (n_405));
  AN21X1 g998(.A (n_394), .B (n_321), .C (n_360), .Q (n_404));
  AN21X1 g999(.A (n_394), .B (n_298), .C (n_336), .Q (n_403));
  AN21X1 g1000(.A (n_394), .B (n_350), .C (n_373), .Q (n_402));
  EN2X1 g1001(.A (n_393), .B (n_270), .Q (out_0[14]));
  EN2X1 g1003(.A (n_389), .B (n_253), .Q (out_0[10]));
  NA2X2 g1005(.A (n_396), .B (n_315), .Q (n_401));
  EN2X1 g1006(.A (n_392), .B (n_271), .Q (out_0[15]));
  EN2X1 g1007(.A (n_391), .B (n_248), .Q (out_0[12]));
  EN2X1 g1008(.A (n_169), .B (n_249), .Q (out_0[13]));
  AN21X1 g1009(.A (n_394), .B (n_352), .C (n_375), .Q (n_400));
  NO2X1 g1010(.A (n_396), .B (n_341), .Q (n_399));
  AN21X1 g1011(.A (n_394), .B (n_353), .C (n_372), .Q (n_398));
  AN21X1 g1012(.A (n_394), .B (n_349), .C (n_376), .Q (n_397));
  NO2X2 g1013(.A (n_395), .B (n_314), .Q (n_396));
  INX8 g1014(.A (n_395), .Q (n_394));
  NO2X4 g1015(.A (n_387), .B (n_366), .Q (n_395));
  AN31X1 g1016(.A (n_275), .B (n_313), .C (n_168), .D (n_367), .Q
       (n_393));
  AO31X1 g1018(.A (n_313), .B (n_316), .C (n_168), .D (n_370), .Q
       (n_392));
  EN2X1 g1019(.A (n_168), .B (n_247), .Q (out_0[8]));
  AO21X1 g1020(.A (n_168), .B (n_313), .C (n_355), .Q (n_391));
  AO321X2 g1021(.A (n_175), .B (n_256), .C (n_168), .D (n_175), .E
       (n_306), .F (n_229), .Q (n_390));
  AN21X1 g1022(.A (n_168), .B (n_256), .C (n_306), .Q (n_389));
  ON21X1 g1023(.A (n_167), .B (n_184), .C (n_183), .Q (n_388));
  NO2X2 g1024(.A (n_167), .B (n_329), .Q (n_387));
  EN2X1 g1025(.A (n_385), .B (n_269), .Q (out_0[6]));
  EN2X1 g1026(.A (n_386), .B (n_268), .Q (out_0[7]));
  EN2X1 g1027(.A (n_383), .B (n_242), .Q (out_0[5]));
  INX2 g1030(.A (n_167), .Q (n_168));
  NO2X4 g1031(.A (n_432), .B (n_440), .Q (n_167));
  AN31X1 g1032(.A (n_260), .B (n_212), .C (n_380), .D (n_335), .Q
       (n_386));
  NO2X1 g1033(.A (n_382), .B (n_303), .Q (n_385));
  AN21X1 g1035(.A (n_380), .B (n_188), .C (n_193), .Q (n_383));
  EN2X1 g1036(.A (n_381), .B (n_244), .Q (out_0[4]));
  NO2X1 g1037(.A (n_381), .B (n_261), .Q (n_382));
  INX2 g1038(.A (n_380), .Q (n_381));
  EO2X1 g1039(.A (n_243), .B (n_371), .Q (out_0[3]));
  NA2X4 g1040(.A (n_379), .B (n_204), .Q (n_380));
  NA2X2 g1041(.A (n_371), .B (n_203), .Q (n_379));
  EN2X0 g1042(.A (n_365), .B (n_95), .Q (out_0[2]));
  ON21X1 g1043(.A (n_364), .B (n_255), .C (n_307), .Q (n_378));
  ON21X1 g1044(.A (n_364), .B (n_173), .C (n_215), .Q (n_377));
  ON21X1 g1045(.A (n_364), .B (n_312), .C (n_344), .Q (n_376));
  ON211X1 g1046(.A (n_364), .B (n_318), .C (n_324), .D (n_223), .Q
       (n_375));
  ON21X1 g1047(.A (n_364), .B (n_333), .C (n_368), .Q (n_374));
  ON21X1 g1048(.A (n_364), .B (n_332), .C (n_369), .Q (n_373));
  ON211X1 g1049(.A (n_364), .B (n_334), .C (n_359), .D (n_227), .Q
       (n_372));
  NO2I1X2 g1050(.B (n_365), .AN (n_95), .Q (n_371));
  ON211X1 g1051(.A (n_305), .B (n_206), .C (n_357), .D (n_224), .Q
       (n_370));
  AN21X1 g1052(.A (n_436), .B (n_276), .C (n_308), .Q (n_369));
  AN21X1 g1053(.A (n_436), .B (n_319), .C (n_348), .Q (n_368));
  AO21X1 g1054(.A (n_355), .B (n_275), .C (n_304), .Q (n_367));
  NA2X4 g1055(.A (n_358), .B (n_435), .Q (n_366));
  INX1 g1056(.A (n_364), .Q (n_363));
  AN21X1 g1057(.A (n_341), .B (n_315), .C (n_340), .Q (n_362));
  ON21X1 g1058(.A (n_437), .B (n_274), .C (n_166), .Q (n_361));
  ON21X1 g1059(.A (n_437), .B (n_177), .C (n_222), .Q (n_360));
  AN21X1 g1061(.A (n_464), .B (n_200), .C (n_201), .Q (n_365));
  NO2X4 g1062(.A (n_356), .B (n_434), .Q (n_364));
  NA2X1 g1063(.A (n_436), .B (n_214), .Q (n_359));
  NA2X2 g1064(.A (n_355), .B (n_317), .Q (n_358));
  NA2X1 g1065(.A (n_355), .B (n_316), .Q (n_357));
  NO2X1 g1066(.A (n_437), .B (n_320), .Q (n_356));
  NO2X1 g1067(.A (n_331), .B (n_173), .Q (n_354));
  NO2X1 g1068(.A (n_334), .B (n_331), .Q (n_353));
  NO2X1 g1069(.A (n_331), .B (n_318), .Q (n_352));
  NO2X1 g1070(.A (n_331), .B (n_255), .Q (n_351));
  NO2X1 g1071(.A (n_332), .B (n_331), .Q (n_350));
  NO2X1 g1072(.A (n_331), .B (n_312), .Q (n_349));
  ON21X1 g1073(.A (n_309), .B (n_228), .C (n_232), .Q (n_348));
  NO2X1 g1074(.A (n_333), .B (n_331), .Q (n_347));
  NA2X4 g1075(.A (n_326), .B (n_297), .Q (n_355));
  INX1 g1077(.A (n_436), .Q (n_344));
  INX1 g1078(.A (n_437), .Q (n_341));
  ON21X1 g1079(.A (n_166), .B (n_210), .C (n_226), .Q (n_340));
  ON21X1 g1084(.A (n_302), .B (n_174), .C (n_185), .Q (n_336));
  AO21X1 g1085(.A (n_303), .B (n_212), .C (n_230), .Q (n_335));
  INX2 g1089(.A (n_330), .Q (n_331));
  NA2X1 g1090(.A (n_317), .B (n_313), .Q (n_329));
  NO2X1 g1091(.A (n_314), .B (n_274), .Q (n_328));
  NA2X1 g1092(.A (n_311), .B (n_214), .Q (n_334));
  NA2X1 g1093(.A (n_311), .B (n_319), .Q (n_333));
  NA2X1 g1094(.A (n_311), .B (n_276), .Q (n_332));
  NO2X2 g1095(.A (n_320), .B (n_314), .Q (n_330));
  NA2X1 g1097(.A (n_306), .B (n_277), .Q (n_326));
  OR2X1 g1099(.A (n_307), .B (n_207), .Q (n_324));
  NO2X1 g1102(.A (n_314), .B (n_177), .Q (n_321));
  INX1 g1103(.A (n_311), .Q (n_312));
  OR2X2 g1105(.A (n_292), .B (n_274), .Q (n_320));
  NO2I1X1 g1106(.B (n_228), .AN (n_276), .Q (n_319));
  OR2X1 g1107(.A (n_255), .B (n_207), .Q (n_318));
  NO2I1X2 g1108(.B (n_296), .AN (n_275), .Q (n_317));
  NO2I1X1 g1109(.B (n_206), .AN (n_275), .Q (n_316));
  NO2X1 g1110(.A (n_274), .B (n_210), .Q (n_315));
  NA2X1 g1111(.A (n_262), .B (n_257), .Q (n_314));
  AND2X4 g1112(.A (n_277), .B (n_256), .Q (n_313));
  NO2X1 g1113(.A (n_295), .B (n_255), .Q (n_311));
  INX1 g1114(.A (n_308), .Q (n_309));
  INX1 g1115(.A (n_305), .Q (n_304));
  INX1 g1116(.A (n_302), .Q (n_301));
  NO2I1X1 g1119(.B (n_174), .AN (n_257), .Q (n_298));
  AN21X1 g1120(.A (n_229), .B (n_195), .C (n_197), .Q (n_297));
  ON21X1 g1121(.A (n_225), .B (n_227), .C (n_236), .Q (n_308));
  OA21X2 g1122(.A (n_186), .B (n_215), .C (n_198), .Q (n_307));
  ON21X1 g1123(.A (n_191), .B (n_183), .C (n_238), .Q (n_306));
  OA21X2 g1125(.A (n_216), .B (n_219), .C (n_233), .Q (n_305));
  ON21X1 g1126(.A (n_189), .B (n_194), .C (n_205), .Q (n_303));
  NO2X2 g1127(.A (n_254), .B (n_199), .Q (n_302));
  OR2X2 g1140(.A (n_206), .B (n_220), .Q (n_296));
  OR2X1 g1141(.A (n_217), .B (n_207), .Q (n_295));
  NO2I1X1 g1142(.B (n_191), .AN (n_238), .Q (n_294));
  NO2I1X1 g1143(.B (n_221), .AN (n_235), .Q (n_293));
  NA2I1X1 g1144(.B (n_234), .AN (n_220), .Q (n_271));
  NO2I1X1 g1145(.B (n_206), .AN (n_224), .Q (n_270));
  OR2X1 g1146(.A (n_210), .B (n_221), .Q (n_292));
  NO2I1X1 g1147(.B (n_210), .AN (n_226), .Q (n_290));
  AND2X1 g1148(.A (n_212), .B (n_231), .Q (n_269));
  NO2X1 g1149(.A (n_192), .B (n_211), .Q (n_288));
  NO2I1X1 g1150(.B (n_207), .AN (n_223), .Q (n_287));
  NO2I1X1 g1151(.B (n_228), .AN (n_232), .Q (n_286));
  NO2I1X1 g1152(.B (n_217), .AN (n_239), .Q (n_284));
  NO2I1X1 g1153(.B (n_190), .AN (n_237), .Q (n_282));
  NO2I1X1 g1154(.B (n_192), .AN (n_202), .Q (n_268));
  NO2I1X1 g1155(.B (n_225), .AN (n_236), .Q (n_280));
  NA2X1 g1156(.A (n_214), .B (n_227), .Q (n_278));
  NO2X1 g1157(.A (n_176), .B (n_196), .Q (n_277));
  NO2X1 g1158(.A (n_213), .B (n_225), .Q (n_276));
  NO2X1 g1159(.A (n_208), .B (n_216), .Q (n_275));
  OR2X2 g1160(.A (n_177), .B (n_182), .Q (n_274));
  INX1 g1164(.A (n_262), .Q (n_263));
  INX1 g1165(.A (n_261), .Q (n_260));
  NO2X1 g1167(.A (n_180), .B (n_187), .Q (n_254));
  NO2X1 g1168(.A (n_229), .B (n_176), .Q (n_253));
  NA2I1X1 g1169(.B (n_185), .AN (n_174), .Q (n_252));
  NA2I1X1 g1170(.B (n_215), .AN (n_173), .Q (n_251));
  NO2I1X1 g1171(.B (n_182), .AN (n_240), .Q (n_266));
  NA2I1X1 g1172(.B (n_222), .AN (n_177), .Q (n_250));
  NA2I1X1 g1173(.B (n_233), .AN (n_216), .Q (n_249));
  NA2X1 g1174(.A (n_209), .B (n_219), .Q (n_248));
  NO2I1X1 g1175(.B (n_186), .AN (n_198), .Q (n_265));
  NO2X1 g1176(.A (n_196), .B (n_197), .Q (n_264));
  NO2X2 g1177(.A (n_190), .B (n_174), .Q (n_262));
  NA2I1X1 g1178(.B (n_183), .AN (n_184), .Q (n_247));
  NO2I1X1 g1179(.B (n_181), .AN (n_179), .Q (n_246));
  NO2I1X1 g1180(.B (n_201), .AN (n_200), .Q (n_245));
  NA2I1X1 g1181(.B (n_188), .AN (n_189), .Q (n_261));
  AND2X1 g1183(.A (n_188), .B (n_194), .Q (n_244));
  AND2X1 g1184(.A (n_203), .B (n_204), .Q (n_243));
  NO2I1X1 g1185(.B (n_189), .AN (n_205), .Q (n_242));
  OR2X1 g1186(.A (n_199), .B (n_187), .Q (n_241));
  NO2X1 g1187(.A (n_178), .B (n_187), .Q (n_257));
  NO2X1 g1188(.A (n_191), .B (n_184), .Q (n_256));
  OR2X1 g1189(.A (n_173), .B (n_186), .Q (n_255));
  INX1 g1190(.A (n_231), .Q (n_230));
  INX1 g1191(.A (n_219), .Q (n_218));
  INX1 g1192(.A (n_213), .Q (n_214));
  INX1 g1193(.A (n_211), .Q (n_212));
  INX1 g1194(.A (n_208), .Q (n_209));
  NA2X1 g1195(.A (n_460), .B (n_148), .Q (n_240));
  NA2X1 g1196(.A (n_442), .B (n_155), .Q (n_239));
  NA2X1 g1197(.A (n_450), .B (n_135), .Q (n_238));
  NA2X1 g1198(.A (n_114), .B (n_146), .Q (n_237));
  NA2X1 g1199(.A (n_444), .B (n_157), .Q (n_236));
  NA2X1 g1200(.A (n_118), .B (n_461), .Q (n_235));
  NA2X1 g1201(.A (n_109), .B (n_142), .Q (n_234));
  NA2X1 g1202(.A (n_456), .B (n_139), .Q (n_233));
  NA2X1 g1203(.A (n_446), .B (n_443), .Q (n_232));
  NA2X1 g1204(.A (n_99), .B (n_447), .Q (n_231));
  AND2X1 g1205(.A (n_452), .B (n_449), .Q (n_229));
  NO2X1 g1206(.A (n_446), .B (n_443), .Q (n_228));
  NA2X1 g1207(.A (n_124), .B (n_441), .Q (n_227));
  NA2X1 g1208(.A (n_462), .B (n_459), .Q (n_226));
  NO2X1 g1209(.A (n_444), .B (n_157), .Q (n_225));
  NA2X1 g1210(.A (n_108), .B (n_455), .Q (n_224));
  NA2X1 g1211(.A (n_121), .B (n_154), .Q (n_223));
  NA2X1 g1212(.A (n_115), .B (n_147), .Q (n_222));
  NO2X1 g1213(.A (n_118), .B (n_461), .Q (n_221));
  NO2X1 g1214(.A (n_109), .B (n_142), .Q (n_220));
  NA2X1 g1215(.A (n_106), .B (n_453), .Q (n_219));
  NO2X1 g1216(.A (n_442), .B (n_155), .Q (n_217));
  NO2X2 g1217(.A (n_456), .B (n_139), .Q (n_216));
  NA2X1 g1218(.A (n_119), .B (n_151), .Q (n_215));
  NO2X1 g1219(.A (n_124), .B (n_441), .Q (n_213));
  NO2X2 g1220(.A (n_99), .B (n_447), .Q (n_211));
  NO2X1 g1221(.A (n_462), .B (n_459), .Q (n_210));
  NO2X1 g1222(.A (n_106), .B (n_453), .Q (n_208));
  NO2X1 g1223(.A (n_121), .B (n_154), .Q (n_207));
  NO2X2 g1224(.A (n_108), .B (n_455), .Q (n_206));
  INX1 g1225(.A (n_196), .Q (n_195));
  INX1 g1226(.A (n_194), .Q (n_193));
  INX1 g1227(.A (n_180), .Q (n_181));
  INX1 g1228(.A (n_178), .Q (n_179));
  INX1 g1229(.A (n_176), .Q (n_175));
  NA2X1 g1233(.A (n_448), .B (n_131), .Q (n_205));
  NA2X1 g1234(.A (n_96), .B (n_128), .Q (n_204));
  OR2X2 g1235(.A (n_96), .B (n_128), .Q (n_203));
  NA2X1 g1236(.A (n_101), .B (n_133), .Q (n_202));
  AND2X1 g1237(.A (in_1[1]), .B (in_0[1]), .Q (n_201));
  OR2X2 g1238(.A (in_1[1]), .B (in_0[1]), .Q (n_200));
  AND2X1 g1239(.A (n_144), .B (n_458), .Q (n_199));
  NA2X1 g1240(.A (n_120), .B (n_153), .Q (n_198));
  AND2X1 g1241(.A (n_454), .B (n_451), .Q (n_197));
  NO2X2 g1242(.A (n_454), .B (n_451), .Q (n_196));
  NA2X1 g1243(.A (n_97), .B (n_129), .Q (n_194));
  NO2X2 g1244(.A (n_101), .B (n_133), .Q (n_192));
  NO2X1 g1245(.A (n_450), .B (n_135), .Q (n_191));
  NO2X2 g1246(.A (n_114), .B (n_146), .Q (n_190));
  NO2X1 g1247(.A (n_448), .B (n_131), .Q (n_189));
  OR2X1 g1248(.A (n_97), .B (n_129), .Q (n_188));
  NO2X2 g1249(.A (n_458), .B (n_144), .Q (n_187));
  NO2X1 g1250(.A (n_120), .B (n_153), .Q (n_186));
  NA2X1 g1251(.A (n_113), .B (n_457), .Q (n_185));
  NO2X1 g1252(.A (n_102), .B (n_134), .Q (n_184));
  NA2X1 g1253(.A (n_102), .B (n_134), .Q (n_183));
  NO2X1 g1254(.A (n_460), .B (n_148), .Q (n_182));
  NA2X1 g1255(.A (n_110), .B (n_143), .Q (n_180));
  NO2X1 g1256(.A (n_110), .B (n_143), .Q (n_178));
  NO2X1 g1257(.A (n_115), .B (n_147), .Q (n_177));
  NO2X1 g1258(.A (n_452), .B (n_449), .Q (n_176));
  NO2X2 g1259(.A (n_113), .B (n_457), .Q (n_174));
  NO2X1 g1260(.A (n_119), .B (n_151), .Q (n_173));
  EO2X1 g300(.A (n_388), .B (n_294), .Q (out_0[9]));
  EN2X1 g1261(.A (n_412), .B (n_293), .Q (out_0[23]));
  EN2X1 g1262(.A (n_407), .B (n_287), .Q (out_0[26]));
  EN2X1 g1263(.A (n_402), .B (n_286), .Q (out_0[30]));
  EN2X1 g1264(.A (n_406), .B (n_265), .Q (out_0[25]));
  EO2X1 g1265(.A (n_390), .B (n_264), .Q (out_0[11]));
  OA21X1 g1267(.A (n_182), .B (n_222), .C (n_240), .Q (n_166));
  AO321X1 g1269(.A (n_209), .B (n_313), .C (n_168), .D (n_209), .E
       (n_355), .F (n_218), .Q (n_169));
  EN2X1 g1280(.A (n_404), .B (n_266), .Q (out_0[21]));
  EO2X1 g1281(.A (n_408), .B (n_438), .Q (out_0[31]));
  EN2X1 g1282(.A (n_398), .B (n_280), .Q (out_0[29]));
  EN2X1 g1283(.A (n_405), .B (n_290), .Q (out_0[22]));
  EO2X1 g1284(.A (n_397), .B (n_278), .Q (out_0[28]));
  EN2X1 g1285(.A (n_400), .B (n_284), .Q (out_0[27]));
  EN2X1 g1286(.A (n_403), .B (n_282), .Q (out_0[19]));
  NO3I1X2 g1288(.B (n_261), .C (n_381), .AN (n_288), .Q (n_432));
  EO2X1 g1289(.A (n_245), .B (n_464), .Q (out_0[1]));
  ON221X1 g1290(.A (n_166), .B (n_292), .C (n_221), .D (n_226), .E
       (n_235), .Q (n_434));
  OA221X2 g1291(.A (n_305), .B (n_296), .C (n_220), .D (n_224), .E
       (n_234), .Q (n_435));
  ON221X1 g1292(.A (n_307), .B (n_295), .C (n_217), .D (n_223), .E
       (n_239), .Q (n_436));
  OA221X4 g1293(.A (n_263), .B (n_302), .C (n_190), .D (n_185), .E
       (n_237), .Q (n_437));
  EN3X1 g1294(.A (in_1[31]), .B (in_0[31]), .C (n_445), .Q (n_438));
  AO21X2 g1295(.A (n_303), .B (n_288), .C (n_439), .Q (n_440));
  ON21X1 g3(.A (n_192), .B (n_231), .C (n_202), .Q (n_439));
  HAX2 g1296(.A (in_1[27]), .B (in_0[27]), .S (n_442), .CO (n_441));
  HAX2 g1297(.A (in_1[29]), .B (in_0[29]), .S (n_444), .CO (n_443));
  HAX2 g1298(.A (in_1[30]), .B (in_0[30]), .S (n_446), .CO (n_445));
  HAX2 g2(.A (in_1[5]), .B (in_0[5]), .S (n_448), .CO (n_447));
  HAX2 g1299(.A (in_1[9]), .B (in_0[9]), .S (n_450), .CO (n_449));
  HAX2 g1300(.A (in_1[10]), .B (in_0[10]), .S (n_452), .CO (n_451));
  HAX2 g1301(.A (in_1[11]), .B (in_0[11]), .S (n_454), .CO (n_453));
  HAX2 g1302(.A (in_1[13]), .B (in_0[13]), .S (n_456), .CO (n_455));
  HAX2 g1303(.A (in_1[17]), .B (in_0[17]), .S (n_458), .CO (n_457));
  HAX2 g1304(.A (in_1[21]), .B (in_0[21]), .S (n_460), .CO (n_459));
  HAX2 g1305(.A (in_1[22]), .B (in_0[22]), .S (n_462), .CO (n_461));
  FAX4 g1306(.A (in_1[0]), .B (in_0[0]), .CI (in_2[0]), .S (out_0[0]),
       .CO (n_464));
endmodule

module rvsteel_core(clock, reset, halt, rw_address, read_data,
     read_request, read_response, write_data, write_strobe,
     write_request, write_response, irq_external,
     irq_external_response, irq_timer, irq_timer_response,
     irq_software, irq_software_response, irq_fast, irq_fast_response,
     real_time_clock);
  input clock, reset, halt, read_response, write_response,
       irq_external, irq_timer, irq_software;
  input [31:0] read_data;
  input [15:0] irq_fast;
  input [63:0] real_time_clock;
  output [31:0] rw_address, write_data;
  output read_request, write_request, irq_external_response,
       irq_timer_response, irq_software_response;
  output [3:0] write_strobe;
  output [15:0] irq_fast_response;
  wire clock, reset, halt, read_response, write_response, irq_external,
       irq_timer, irq_software;
  wire [31:0] read_data;
  wire [15:0] irq_fast;
  wire [63:0] real_time_clock;
  wire [31:0] rw_address, write_data;
  wire read_request, write_request, irq_external_response,
       irq_timer_response, irq_software_response;
  wire [3:0] write_strobe;
  wire [15:0] irq_fast_response;
  wire [31:0] alu_sra_result;
  wire [31:0] prev_rw_address;
  wire [31:0] csr_mscratch;
  wire [31:0] prev_instruction;
  wire [3:0] current_state;
  wire [31:0] instruction;
  wire [63:0] csr_utime;
  wire [31:0] csr_data_out;
  wire [31:0] prev_instruction_address;
  wire [31:0] csr_mtval;
  wire [31:0] csr_mcause;
  wire [3:0] prev_write_strobe;
  wire [31:0] program_counter;
  wire [31:0] alu_2nd_operand;
  wire [31:0] prev_write_data;
  wire [31:0] csr_mtvec;
  wire [63:0] csr_mcycle;
  wire [63:0] csr_minstret;
  wire [4:0] csr_mcause_code;
  wire UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2,
       UNCONNECTED3, UNCONNECTED4, UNCONNECTED5, UNCONNECTED6;
  wire UNCONNECTED7, UNCONNECTED8, UNCONNECTED9, UNCONNECTED10,
       UNCONNECTED11, UNCONNECTED12, UNCONNECTED13, UNCONNECTED14;
  wire UNCONNECTED15, UNCONNECTED16, UNCONNECTED17, UNCONNECTED18,
       UNCONNECTED19, UNCONNECTED20, UNCONNECTED21, UNCONNECTED22;
  wire UNCONNECTED23, UNCONNECTED24, UNCONNECTED25, UNCONNECTED_HIER_Z,
       UNCONNECTED_HIER_Z0, UNCONNECTED_HIER_Z1, UNCONNECTED_HIER_Z2,
       UNCONNECTED_HIER_Z3;
  wire UNCONNECTED_HIER_Z4, UNCONNECTED_HIER_Z5, UNCONNECTED_HIER_Z6,
       UNCONNECTED_HIER_Z7, UNCONNECTED_HIER_Z8, UNCONNECTED_HIER_Z9,
       UNCONNECTED_HIER_Z10, UNCONNECTED_HIER_Z11;
  wire UNCONNECTED_HIER_Z12, UNCONNECTED_HIER_Z13,
       UNCONNECTED_HIER_Z14, UNCONNECTED_HIER_Z15,
       UNCONNECTED_HIER_Z16, UNCONNECTED_HIER_Z17,
       UNCONNECTED_HIER_Z18, UNCONNECTED_HIER_Z19;
  wire UNCONNECTED_HIER_Z20, UNCONNECTED_HIER_Z21,
       UNCONNECTED_HIER_Z22, UNCONNECTED_HIER_Z23,
       UNCONNECTED_HIER_Z24, UNCONNECTED_HIER_Z25,
       UNCONNECTED_HIER_Z26, UNCONNECTED_HIER_Z27;
  wire UNCONNECTED_HIER_Z28, UNCONNECTED_HIER_Z29,
       UNCONNECTED_HIER_Z30, UNCONNECTED_HIER_Z31,
       UNCONNECTED_HIER_Z32, UNCONNECTED_HIER_Z33, add_459_21_n_642,
       add_459_21_n_645;
  wire add_459_21_n_648, add_459_21_n_652, add_459_21_n_654,
       add_459_21_n_658, add_459_21_n_660, add_459_21_n_662,
       add_459_21_n_664, add_459_21_n_666;
  wire add_459_21_n_668, add_459_21_n_670, add_459_21_n_672,
       add_459_21_n_674, add_459_21_n_676, add_459_21_n_677,
       add_459_21_n_682, add_459_21_n_684;
  wire add_459_21_n_685, add_459_21_n_692, add_459_21_n_693,
       add_459_21_n_700, add_459_21_n_701, add_459_21_n_708,
       add_459_21_n_709, add_459_21_n_715;
  wire add_459_21_n_721, add_459_21_n_727, add_463_14_n_597,
       add_463_14_n_599, add_463_14_n_600, add_463_14_n_601,
       add_463_14_n_603, add_463_14_n_605;
  wire add_463_14_n_606, add_463_14_n_607, add_463_14_n_609,
       add_463_14_n_610, add_463_14_n_618, add_463_14_n_619,
       add_463_14_n_620, add_463_14_n_622;
  wire add_463_14_n_623, add_463_14_n_625, add_463_14_n_628,
       add_463_14_n_632, add_463_14_n_634, add_463_14_n_636,
       add_463_14_n_639, add_463_14_n_640;
  wire add_463_14_n_641, add_463_14_n_646, add_463_14_n_647,
       add_463_14_n_648, add_463_14_n_649, add_463_14_n_653,
       add_463_14_n_655, add_463_14_n_656;
  wire add_463_14_n_659, add_463_14_n_660, add_463_14_n_662,
       add_463_14_n_663, add_463_14_n_664, add_463_14_n_666,
       add_463_14_n_667, add_463_14_n_672;
  wire add_463_14_n_673, add_463_14_n_675, add_463_14_n_676,
       add_463_14_n_678, add_463_14_n_680, add_463_14_n_681,
       add_463_14_n_682, add_463_14_n_683;
  wire add_463_14_n_684, add_463_14_n_688, add_463_14_n_691,
       add_463_14_n_693, add_463_14_n_695, add_463_14_n_697,
       add_463_14_n_698, add_463_14_n_699;
  wire add_463_14_n_701, add_463_14_n_702, add_463_14_n_703,
       add_463_14_n_705, add_463_14_n_708, add_463_14_n_709,
       add_463_14_n_710, add_463_14_n_711;
  wire add_463_14_n_714, add_463_14_n_717, add_463_14_n_720,
       add_463_14_n_721, add_463_14_n_722, add_463_14_n_723,
       add_463_14_n_724, add_463_14_n_725;
  wire add_463_14_n_726, add_463_14_n_730, add_463_14_n_740,
       add_463_14_n_741, add_463_14_n_746, add_463_14_n_748,
       add_463_14_n_749, add_463_14_n_750;
  wire add_463_14_n_751, add_463_14_n_752, add_463_14_n_753,
       add_463_14_n_754, add_463_14_n_755, add_463_14_n_756,
       add_463_14_n_757, add_463_14_n_758;
  wire add_463_14_n_759, add_463_14_n_760, add_463_14_n_761,
       add_463_14_n_762, add_463_14_n_763, add_463_14_n_764,
       add_463_14_n_776, add_463_14_n_777;
  wire add_463_14_n_778, add_463_14_n_779, add_463_14_n_780,
       add_463_14_n_781, add_463_14_n_782, add_463_14_n_783,
       add_463_14_n_784, add_463_14_n_785;
  wire add_463_14_n_792, add_463_14_n_793, add_463_14_n_794,
       add_463_14_n_795, add_463_14_n_796, add_463_14_n_797,
       add_463_14_n_798, add_463_14_n_799;
  wire add_463_14_n_800, add_463_14_n_801, add_463_14_n_802,
       add_463_14_n_804, add_463_14_n_807, add_463_14_n_810,
       add_463_14_n_811, add_463_14_n_812;
  wire add_463_14_n_813, add_463_14_n_814, add_463_14_n_817,
       add_463_14_n_821, add_463_14_n_823, add_463_14_n_826,
       add_463_14_n_828, add_463_14_n_836;
  wire add_463_14_n_837, add_463_14_n_838, add_463_14_n_839,
       add_463_14_n_840, add_463_14_n_843, add_463_14_n_845,
       add_463_14_n_847, add_463_14_n_850;
  wire add_463_14_n_853, add_463_14_n_855, add_463_14_n_857,
       add_463_14_n_859, add_463_14_n_862, add_463_14_n_864,
       add_463_14_n_866, add_463_14_n_868;
  wire add_463_14_n_870, add_463_14_n_872, add_463_14_n_875,
       add_463_14_n_877, add_463_14_n_880, add_463_14_n_883,
       add_463_14_n_884, add_463_14_n_885;
  wire add_463_14_n_886, add_463_14_n_887, add_463_14_n_888,
       add_463_14_n_889, add_463_14_n_890, add_463_14_n_891,
       add_463_14_n_892, add_463_14_n_893;
  wire add_463_14_n_894, add_463_14_n_895, add_463_14_n_896,
       add_463_14_n_897, add_463_14_n_898, add_463_14_n_899,
       add_463_14_n_900, add_463_14_n_901;
  wire add_463_14_n_902, add_463_14_n_903, add_463_14_n_904,
       add_463_14_n_905, add_463_14_n_906, add_463_14_n_907,
       add_463_14_n_908, add_463_14_n_909;
  wire add_463_14_n_910, add_463_14_n_911, add_463_14_n_912,
       add_463_14_n_913, add_463_14_n_914, add_463_14_n_915,
       add_463_14_n_916, add_463_14_n_917;
  wire add_463_14_n_936, add_463_14_n_937, add_463_14_n_938,
       add_463_14_n_940, add_463_14_n_941, add_463_14_n_942,
       add_463_14_n_943, add_463_14_n_944;
  wire add_463_14_n_945, add_463_14_n_946, add_463_14_n_947,
       add_463_14_n_948, add_463_14_n_949, add_463_14_n_950,
       add_463_14_n_951, add_463_14_n_952;
  wire add_463_14_n_953, add_463_14_n_954, add_463_14_n_955,
       add_463_14_n_956, add_463_14_n_957, add_463_14_n_958,
       add_463_14_n_959, add_463_14_n_960;
  wire add_463_14_n_961, add_463_14_n_962, add_463_14_n_963,
       add_463_14_n_964, add_463_14_n_965, add_463_14_n_966,
       add_463_14_n_967, add_463_14_n_968;
  wire add_463_14_n_969, add_463_14_n_970, add_463_14_n_971,
       add_463_14_n_972, add_463_14_n_973, add_463_14_n_974,
       add_463_14_n_1078, add_464_21_n_596;
  wire add_464_21_n_597, add_464_21_n_599, add_464_21_n_600,
       add_464_21_n_602, add_464_21_n_605, add_464_21_n_608,
       add_464_21_n_611, add_464_21_n_621;
  wire add_464_21_n_622, add_464_21_n_625, add_464_21_n_626,
       add_464_21_n_627, add_464_21_n_632, add_464_21_n_634,
       add_464_21_n_637, add_464_21_n_638;
  wire add_464_21_n_639, add_464_21_n_642, add_464_21_n_643,
       add_464_21_n_645, add_464_21_n_648, add_464_21_n_653,
       add_464_21_n_654, add_464_21_n_655;
  wire add_464_21_n_657, add_464_21_n_661, add_464_21_n_664,
       add_464_21_n_665, add_464_21_n_667, add_464_21_n_669,
       add_464_21_n_674, add_464_21_n_676;
  wire add_464_21_n_678, add_464_21_n_679, add_464_21_n_680,
       add_464_21_n_685, add_464_21_n_686, add_464_21_n_687,
       add_464_21_n_690, add_464_21_n_691;
  wire add_464_21_n_693, add_464_21_n_695, add_464_21_n_697,
       add_464_21_n_701, add_464_21_n_702, add_464_21_n_703,
       add_464_21_n_704, add_464_21_n_706;
  wire add_464_21_n_708, add_464_21_n_713, add_464_21_n_714,
       add_464_21_n_717, add_464_21_n_720, add_464_21_n_721,
       add_464_21_n_723, add_464_21_n_725;
  wire add_464_21_n_726, add_464_21_n_727, add_464_21_n_728,
       add_464_21_n_729, add_464_21_n_730, add_464_21_n_731,
       add_464_21_n_733, add_464_21_n_734;
  wire add_464_21_n_736, add_464_21_n_737, add_464_21_n_738,
       add_464_21_n_745, add_464_21_n_746, add_464_21_n_747,
       add_464_21_n_748, add_464_21_n_749;
  wire add_464_21_n_750, add_464_21_n_751, add_464_21_n_752,
       add_464_21_n_753, add_464_21_n_754, add_464_21_n_755,
       add_464_21_n_756, add_464_21_n_757;
  wire add_464_21_n_765, add_464_21_n_766, add_464_21_n_767,
       add_464_21_n_768, add_464_21_n_769, add_464_21_n_770,
       add_464_21_n_771, add_464_21_n_772;
  wire add_464_21_n_775, add_464_21_n_777, add_464_21_n_779,
       add_464_21_n_782, add_464_21_n_785, add_464_21_n_788,
       add_464_21_n_790, add_464_21_n_791;
  wire add_464_21_n_793, add_464_21_n_795, add_464_21_n_798,
       add_464_21_n_801, add_464_21_n_804, add_464_21_n_807,
       add_464_21_n_808, add_464_21_n_809;
  wire add_464_21_n_810, add_464_21_n_811, add_464_21_n_812,
       add_464_21_n_813, add_464_21_n_815, add_464_21_n_818,
       add_464_21_n_821, add_464_21_n_823;
  wire add_464_21_n_825, add_464_21_n_827, add_464_21_n_829,
       add_464_21_n_830, add_464_21_n_832, add_464_21_n_835,
       add_464_21_n_838, add_464_21_n_841;
  wire add_464_21_n_844, add_464_21_n_846, add_464_21_n_848,
       add_464_21_n_849, add_464_21_n_850, add_464_21_n_851,
       add_464_21_n_852, add_464_21_n_853;
  wire add_464_21_n_854, add_464_21_n_855, add_464_21_n_856,
       add_464_21_n_857, add_464_21_n_858, add_464_21_n_859,
       add_464_21_n_860, add_464_21_n_861;
  wire add_464_21_n_862, add_464_21_n_863, add_464_21_n_864,
       add_464_21_n_865, add_464_21_n_866, add_464_21_n_867,
       add_464_21_n_868, add_464_21_n_869;
  wire add_464_21_n_870, add_464_21_n_871, add_464_21_n_872,
       add_464_21_n_873, add_464_21_n_874, add_464_21_n_875,
       add_464_21_n_876, add_464_21_n_877;
  wire add_464_21_n_878, add_464_21_n_879, add_464_21_n_880,
       add_464_21_n_881, add_464_21_n_882, add_464_21_n_911,
       add_464_21_n_912, add_464_21_n_913;
  wire add_464_21_n_914, add_464_21_n_915, add_464_21_n_916,
       add_464_21_n_917, add_464_21_n_918, add_464_21_n_919,
       add_464_21_n_920, add_464_21_n_921;
  wire add_464_21_n_922, add_464_21_n_923, add_464_21_n_924,
       add_464_21_n_925, add_464_21_n_926, add_464_21_n_927,
       add_464_21_n_928, add_464_21_n_929;
  wire add_464_21_n_930, add_464_21_n_931, add_464_21_n_932,
       add_464_21_n_933, add_464_21_n_934, add_464_21_n_935,
       add_464_21_n_936, add_464_21_n_937;
  wire add_464_21_n_938, add_464_21_n_939, add_464_21_n_940,
       add_464_21_n_941, add_464_21_n_942, add_464_21_n_943,
       add_464_21_n_944, add_464_21_n_945;
  wire add_464_21_n_946, add_464_21_n_947, add_464_21_n_948,
       add_464_21_n_949, add_1545_30_n_811, add_1545_30_n_814,
       add_1545_30_n_816, add_1545_30_n_821;
  wire add_1545_30_n_825, add_1545_30_n_827, add_1545_30_n_829,
       add_1545_30_n_831, add_1545_30_n_833, add_1545_30_n_835,
       add_1545_30_n_837, add_1545_30_n_840;
  wire add_1545_30_n_843, add_1545_30_n_844, add_1545_30_n_847,
       add_1545_30_n_848, add_1545_30_n_851, add_1545_30_n_854,
       add_1545_30_n_855, add_1545_30_n_858;
  wire add_1545_30_n_860, add_1545_30_n_861, add_1545_30_n_867,
       add_1545_30_n_873, add_1545_30_n_876, add_1545_30_n_878,
       add_1545_30_n_880, add_1545_30_n_882;
  wire add_1545_30_n_883, add_1545_30_n_888, add_1545_30_n_892,
       add_1545_30_n_898, add_1545_30_n_901, add_1545_30_n_904,
       alu_operation_code_39112, branch_type;
  wire csr_mcause_interrupt_flag, flush_37557,
       inc_ADD_UNS_OP5491_6_n_2351, inc_ADD_UNS_OP5491_6_n_2356,
       inc_ADD_UNS_OP5491_6_n_2362, inc_ADD_UNS_OP5491_6_n_2366,
       inc_ADD_UNS_OP5491_6_n_2372, inc_ADD_UNS_OP5491_6_n_2380;
  wire inc_ADD_UNS_OP5491_6_n_2388, inc_ADD_UNS_OP5491_6_n_2393,
       inc_ADD_UNS_OP5491_6_n_2399, inc_ADD_UNS_OP5491_6_n_2401,
       inc_ADD_UNS_OP5491_6_n_2410, inc_ADD_UNS_OP5491_6_n_2419,
       inc_ADD_UNS_OP5491_6_n_2421, inc_ADD_UNS_OP5491_6_n_2424;
  wire inc_ADD_UNS_OP5491_6_n_2431, inc_ADD_UNS_OP5491_6_n_2438,
       inc_ADD_UNS_OP5491_6_n_2440, inc_ADD_UNS_OP5491_6_n_2443,
       inc_ADD_UNS_OP5491_6_n_2446, inc_ADD_UNS_OP5491_6_n_2450,
       inc_ADD_UNS_OP5491_6_n_2452, inc_ADD_UNS_OP5491_6_n_2455;
  wire inc_ADD_UNS_OP5491_6_n_2458, inc_ADD_UNS_OP5491_6_n_2460,
       inc_ADD_UNS_OP5491_6_n_2463, inc_ADD_UNS_OP5491_6_n_2468,
       inc_ADD_UNS_OP5491_6_n_2473, inc_ADD_UNS_OP5491_6_n_2476,
       inc_ADD_UNS_OP5491_6_n_2479, inc_ADD_UNS_OP5491_6_n_2481;
  wire inc_ADD_UNS_OP5491_6_n_2484, inc_ADD_UNS_OP5491_6_n_2489,
       inc_ADD_UNS_OP5491_6_n_2493, inc_ADD_UNS_OP5491_6_n_2497,
       inc_ADD_UNS_OP5491_6_n_2503, inc_ADD_UNS_OP5491_6_n_2507,
       inc_ADD_UNS_OP5491_6_n_2515, inc_ADD_UNS_OP5491_6_n_2517;
  wire inc_ADD_UNS_OP5491_6_n_2521, inc_ADD_UNS_OP5491_6_n_2523,
       inc_ADD_UNS_OP5491_6_n_2526, inc_ADD_UNS_OP5491_6_n_2527,
       inc_ADD_UNS_OP5491_6_n_2531, inc_ADD_UNS_OP5491_6_n_2534,
       inc_ADD_UNS_OP5491_6_n_2537, inc_ADD_UNS_OP5491_6_n_2540;
  wire inc_ADD_UNS_OP5491_6_n_2543, inc_ADD_UNS_OP5491_6_n_2546,
       inc_ADD_UNS_OP5491_6_n_2548, inc_ADD_UNS_OP5491_6_n_2551,
       inc_ADD_UNS_OP5491_6_n_2556, inc_ADD_UNS_OP5491_6_n_2561,
       inc_ADD_UNS_OP5491_6_n_2566, inc_ADD_UNS_OP5491_6_n_2571;
  wire inc_ADD_UNS_OP5491_6_n_2576, inc_ADD_UNS_OP5491_6_n_2581,
       inc_ADD_UNS_OP5491_6_n_2586, inc_ADD_UNS_OP5491_6_n_2591,
       inc_ADD_UNS_OP5491_6_n_2596, inc_ADD_UNS_OP5491_6_n_2601,
       inc_ADD_UNS_OP5491_6_n_2606, inc_ADD_UNS_OP5491_6_n_2611;
  wire inc_ADD_UNS_OP5491_6_n_2615, inc_ADD_UNS_OP5491_6_n_2616,
       inc_ADD_UNS_OP5491_6_n_2620, inc_ADD_UNS_OP5491_6_n_2622,
       inc_ADD_UNS_OP5491_6_n_2625, inc_ADD_UNS_OP5491_6_n_2626,
       inc_ADD_UNS_OP5491_6_n_2628, inc_ADD_UNS_OP5491_6_n_2633;
  wire inc_ADD_UNS_OP5491_6_n_2636, inc_ADD_UNS_OP5491_6_n_2641,
       inc_ADD_UNS_OP5491_6_n_2657, inc_ADD_UNS_OP5491_6_n_2669,
       inc_ADD_UNS_OP5491_6_n_2675, inc_ADD_UNS_OP5491_6_n_2724,
       inc_ADD_UNS_OP5491_6_n_2725, inc_ADD_UNS_OP5492_3_n_2334;
  wire inc_ADD_UNS_OP5492_3_n_2339, inc_ADD_UNS_OP5492_3_n_2344,
       inc_ADD_UNS_OP5492_3_n_2350, inc_ADD_UNS_OP5492_3_n_2356,
       inc_ADD_UNS_OP5492_3_n_2361, inc_ADD_UNS_OP5492_3_n_2366,
       inc_ADD_UNS_OP5492_3_n_2371, inc_ADD_UNS_OP5492_3_n_2377;
  wire inc_ADD_UNS_OP5492_3_n_2380, inc_ADD_UNS_OP5492_3_n_2383,
       inc_ADD_UNS_OP5492_3_n_2388, inc_ADD_UNS_OP5492_3_n_2394,
       inc_ADD_UNS_OP5492_3_n_2399, inc_ADD_UNS_OP5492_3_n_2404,
       inc_ADD_UNS_OP5492_3_n_2409, inc_ADD_UNS_OP5492_3_n_2413;
  wire inc_ADD_UNS_OP5492_3_n_2419, inc_ADD_UNS_OP5492_3_n_2427,
       inc_ADD_UNS_OP5492_3_n_2430, inc_ADD_UNS_OP5492_3_n_2431,
       inc_ADD_UNS_OP5492_3_n_2439, inc_ADD_UNS_OP5492_3_n_2444,
       inc_ADD_UNS_OP5492_3_n_2448, inc_ADD_UNS_OP5492_3_n_2450;
  wire inc_ADD_UNS_OP5492_3_n_2455, inc_ADD_UNS_OP5492_3_n_2459,
       inc_ADD_UNS_OP5492_3_n_2462, inc_ADD_UNS_OP5492_3_n_2465,
       inc_ADD_UNS_OP5492_3_n_2468, inc_ADD_UNS_OP5492_3_n_2472,
       inc_ADD_UNS_OP5492_3_n_2474, inc_ADD_UNS_OP5492_3_n_2476;
  wire inc_ADD_UNS_OP5492_3_n_2479, inc_ADD_UNS_OP5492_3_n_2480,
       inc_ADD_UNS_OP5492_3_n_2485, inc_ADD_UNS_OP5492_3_n_2488,
       inc_ADD_UNS_OP5492_3_n_2490, inc_ADD_UNS_OP5492_3_n_2493,
       inc_ADD_UNS_OP5492_3_n_2497, inc_ADD_UNS_OP5492_3_n_2498;
  wire inc_ADD_UNS_OP5492_3_n_2501, inc_ADD_UNS_OP5492_3_n_2504,
       inc_ADD_UNS_OP5492_3_n_2507, inc_ADD_UNS_OP5492_3_n_2509,
       inc_ADD_UNS_OP5492_3_n_2512, inc_ADD_UNS_OP5492_3_n_2515,
       inc_ADD_UNS_OP5492_3_n_2518, inc_ADD_UNS_OP5492_3_n_2521;
  wire inc_ADD_UNS_OP5492_3_n_2523, inc_ADD_UNS_OP5492_3_n_2533,
       inc_ADD_UNS_OP5492_3_n_2536, inc_ADD_UNS_OP5492_3_n_2539,
       inc_ADD_UNS_OP5492_3_n_2542, inc_ADD_UNS_OP5492_3_n_2545,
       inc_ADD_UNS_OP5492_3_n_2551, inc_ADD_UNS_OP5492_3_n_2553;
  wire inc_ADD_UNS_OP5492_3_n_2556, inc_ADD_UNS_OP5492_3_n_2567,
       inc_ADD_UNS_OP5492_3_n_2571, inc_ADD_UNS_OP5492_3_n_2574,
       inc_ADD_UNS_OP5492_3_n_2580, inc_ADD_UNS_OP5492_3_n_2585,
       inc_ADD_UNS_OP5492_3_n_2608, inc_ADD_UNS_OP5492_3_n_2613;
  wire inc_ADD_UNS_OP5492_3_n_2615, inc_ADD_UNS_OP5492_3_n_2647,
       inc_ADD_UNS_OP5492_3_n_2649, inc_ADD_UNS_OP5492_3_n_2656,
       inc_ADD_UNS_OP5492_3_n_2675, inc_ADD_UNS_OP5492_3_n_2676,
       inc_ADD_UNS_OP_5_n_3370, inc_ADD_UNS_OP_5_n_3387;
  wire inc_ADD_UNS_OP_5_n_3392, inc_ADD_UNS_OP_5_n_3400,
       inc_ADD_UNS_OP_5_n_3411, inc_ADD_UNS_OP_5_n_3415,
       inc_ADD_UNS_OP_5_n_3421, inc_ADD_UNS_OP_5_n_3424,
       inc_ADD_UNS_OP_5_n_3430, inc_ADD_UNS_OP_5_n_3432;
  wire inc_ADD_UNS_OP_5_n_3435, inc_ADD_UNS_OP_5_n_3438,
       inc_ADD_UNS_OP_5_n_3445, inc_ADD_UNS_OP_5_n_3447,
       inc_ADD_UNS_OP_5_n_3453, inc_ADD_UNS_OP_5_n_3463,
       inc_ADD_UNS_OP_5_n_3469, inc_ADD_UNS_OP_5_n_3470;
  wire inc_ADD_UNS_OP_5_n_3474, inc_ADD_UNS_OP_5_n_3476,
       inc_ADD_UNS_OP_5_n_3482, inc_ADD_UNS_OP_5_n_3490,
       inc_ADD_UNS_OP_5_n_3494, inc_ADD_UNS_OP_5_n_3499,
       inc_ADD_UNS_OP_5_n_3505, inc_ADD_UNS_OP_5_n_3509;
  wire inc_ADD_UNS_OP_5_n_3515, inc_ADD_UNS_OP_5_n_3522,
       inc_ADD_UNS_OP_5_n_3527, inc_ADD_UNS_OP_5_n_3530,
       inc_ADD_UNS_OP_5_n_3531, inc_ADD_UNS_OP_5_n_3536,
       inc_ADD_UNS_OP_5_n_3538, inc_ADD_UNS_OP_5_n_3541;
  wire inc_ADD_UNS_OP_5_n_3556, inc_ADD_UNS_OP_5_n_3559,
       inc_ADD_UNS_OP_5_n_3567, inc_ADD_UNS_OP_5_n_3573,
       inc_ADD_UNS_OP_5_n_3574, inc_ADD_UNS_OP_5_n_3580,
       inc_ADD_UNS_OP_5_n_3581, inc_ADD_UNS_OP_5_n_3583;
  wire inc_ADD_UNS_OP_5_n_3590, inc_ADD_UNS_OP_5_n_3597,
       inc_ADD_UNS_OP_5_n_3605, inc_ADD_UNS_OP_5_n_3606,
       inc_ADD_UNS_OP_5_n_3611, inc_ADD_UNS_OP_5_n_3614,
       inc_ADD_UNS_OP_5_n_3616, inc_ADD_UNS_OP_5_n_3621;
  wire inc_ADD_UNS_OP_5_n_3622, inc_ADD_UNS_OP_5_n_3628,
       inc_ADD_UNS_OP_5_n_3631, inc_ADD_UNS_OP_5_n_3637,
       inc_ADD_UNS_OP_5_n_3641, inc_ADD_UNS_OP_5_n_3643,
       inc_ADD_UNS_OP_5_n_3645, inc_ADD_UNS_OP_5_n_3648;
  wire inc_ADD_UNS_OP_5_n_3651, inc_ADD_UNS_OP_5_n_3655,
       inc_ADD_UNS_OP_5_n_3658, inc_ADD_UNS_OP_5_n_3663,
       inc_ADD_UNS_OP_5_n_3664, inc_ADD_UNS_OP_5_n_3665,
       inc_ADD_UNS_OP_5_n_3668, inc_ADD_UNS_OP_5_n_3670;
  wire inc_ADD_UNS_OP_5_n_3676, inc_ADD_UNS_OP_5_n_3681,
       inc_ADD_UNS_OP_5_n_3684, inc_ADD_UNS_OP_5_n_3686,
       inc_ADD_UNS_OP_5_n_3692, inc_ADD_UNS_OP_5_n_3695,
       inc_ADD_UNS_OP_5_n_3697, inc_ADD_UNS_OP_5_n_3701;
  wire inc_ADD_UNS_OP_5_n_3703, inc_ADD_UNS_OP_5_n_3704,
       inc_ADD_UNS_OP_5_n_3708, inc_ADD_UNS_OP_5_n_3711,
       inc_ADD_UNS_OP_5_n_3714, inc_ADD_UNS_OP_5_n_3717,
       inc_ADD_UNS_OP_5_n_3721, inc_ADD_UNS_OP_5_n_3724;
  wire inc_ADD_UNS_OP_5_n_3726, inc_ADD_UNS_OP_5_n_3733,
       inc_ADD_UNS_OP_5_n_3735, inc_ADD_UNS_OP_5_n_3742,
       inc_ADD_UNS_OP_5_n_3746, inc_ADD_UNS_OP_5_n_3748,
       inc_ADD_UNS_OP_5_n_3750, inc_ADD_UNS_OP_5_n_3752;
  wire inc_ADD_UNS_OP_5_n_3756, inc_ADD_UNS_OP_5_n_3760,
       inc_ADD_UNS_OP_5_n_3766, inc_ADD_UNS_OP_5_n_3768,
       inc_ADD_UNS_OP_5_n_3775, inc_ADD_UNS_OP_5_n_3782,
       inc_ADD_UNS_OP_5_n_3785, inc_ADD_UNS_OP_5_n_3789;
  wire inc_ADD_UNS_OP_5_n_3791, inc_ADD_UNS_OP_5_n_3792,
       inc_ADD_UNS_OP_5_n_3793, inc_ADD_UNS_OP_5_n_3795,
       inc_ADD_UNS_OP_5_n_3798, inc_ADD_UNS_OP_5_n_3800,
       inc_ADD_UNS_OP_5_n_3803, inc_ADD_UNS_OP_5_n_3808;
  wire inc_ADD_UNS_OP_5_n_3812, inc_ADD_UNS_OP_5_n_3815,
       inc_ADD_UNS_OP_5_n_3824, inc_ADD_UNS_OP_5_n_3826,
       inc_ADD_UNS_OP_5_n_3832, inc_ADD_UNS_OP_5_n_3834,
       inc_ADD_UNS_OP_5_n_3838, inc_add_1343_59_4_n_3386;
  wire inc_add_1343_59_4_n_3391, inc_add_1343_59_4_n_3403,
       inc_add_1343_59_4_n_3413, inc_add_1343_59_4_n_3419,
       inc_add_1343_59_4_n_3423, inc_add_1343_59_4_n_3428,
       inc_add_1343_59_4_n_3432, inc_add_1343_59_4_n_3435;
  wire inc_add_1343_59_4_n_3440, inc_add_1343_59_4_n_3443,
       inc_add_1343_59_4_n_3446, inc_add_1343_59_4_n_3451,
       inc_add_1343_59_4_n_3457, inc_add_1343_59_4_n_3462,
       inc_add_1343_59_4_n_3468, inc_add_1343_59_4_n_3475;
  wire inc_add_1343_59_4_n_3479, inc_add_1343_59_4_n_3481,
       inc_add_1343_59_4_n_3486, inc_add_1343_59_4_n_3492,
       inc_add_1343_59_4_n_3496, inc_add_1343_59_4_n_3501,
       inc_add_1343_59_4_n_3505, inc_add_1343_59_4_n_3508;
  wire inc_add_1343_59_4_n_3512, inc_add_1343_59_4_n_3519,
       inc_add_1343_59_4_n_3524, inc_add_1343_59_4_n_3527,
       inc_add_1343_59_4_n_3533, inc_add_1343_59_4_n_3536,
       inc_add_1343_59_4_n_3539, inc_add_1343_59_4_n_3544;
  wire inc_add_1343_59_4_n_3551, inc_add_1343_59_4_n_3555,
       inc_add_1343_59_4_n_3558, inc_add_1343_59_4_n_3561,
       inc_add_1343_59_4_n_3572, inc_add_1343_59_4_n_3576,
       inc_add_1343_59_4_n_3578, inc_add_1343_59_4_n_3583;
  wire inc_add_1343_59_4_n_3586, inc_add_1343_59_4_n_3592,
       inc_add_1343_59_4_n_3594, inc_add_1343_59_4_n_3602,
       inc_add_1343_59_4_n_3605, inc_add_1343_59_4_n_3611,
       inc_add_1343_59_4_n_3614, inc_add_1343_59_4_n_3620;
  wire inc_add_1343_59_4_n_3621, inc_add_1343_59_4_n_3624,
       inc_add_1343_59_4_n_3628, inc_add_1343_59_4_n_3629,
       inc_add_1343_59_4_n_3633, inc_add_1343_59_4_n_3635,
       inc_add_1343_59_4_n_3640, inc_add_1343_59_4_n_3642;
  wire inc_add_1343_59_4_n_3646, inc_add_1343_59_4_n_3648,
       inc_add_1343_59_4_n_3649, inc_add_1343_59_4_n_3653,
       inc_add_1343_59_4_n_3656, inc_add_1343_59_4_n_3658,
       inc_add_1343_59_4_n_3660, inc_add_1343_59_4_n_3663;
  wire inc_add_1343_59_4_n_3664, inc_add_1343_59_4_n_3665,
       inc_add_1343_59_4_n_3669, inc_add_1343_59_4_n_3674,
       inc_add_1343_59_4_n_3677, inc_add_1343_59_4_n_3680,
       inc_add_1343_59_4_n_3681, inc_add_1343_59_4_n_3684;
  wire inc_add_1343_59_4_n_3687, inc_add_1343_59_4_n_3693,
       inc_add_1343_59_4_n_3696, inc_add_1343_59_4_n_3718,
       inc_add_1343_59_4_n_3727, inc_add_1343_59_4_n_3736,
       inc_add_1343_59_4_n_3749, inc_add_1343_59_4_n_3758;
  wire inc_add_1343_59_4_n_3766, inc_add_1343_59_4_n_3769,
       inc_add_1343_59_4_n_3775, inc_add_1343_59_4_n_3779,
       inc_add_1343_59_4_n_3784, inc_add_1343_59_4_n_3786,
       inc_add_1343_59_4_n_3788, inc_add_1343_59_4_n_3805;
  wire inc_add_1343_59_4_n_3806, inc_add_1343_59_4_n_3812,
       inc_add_1345_58_1_n_3147, inc_add_1345_58_1_n_3151,
       inc_add_1345_58_1_n_3155, inc_add_1345_58_1_n_3159,
       inc_add_1345_58_1_n_3166, inc_add_1345_58_1_n_3169;
  wire inc_add_1345_58_1_n_3172, inc_add_1345_58_1_n_3175,
       inc_add_1345_58_1_n_3180, inc_add_1345_58_1_n_3185,
       inc_add_1345_58_1_n_3190, inc_add_1345_58_1_n_3195,
       inc_add_1345_58_1_n_3199, inc_add_1345_58_1_n_3202;
  wire inc_add_1345_58_1_n_3205, inc_add_1345_58_1_n_3207,
       inc_add_1345_58_1_n_3210, inc_add_1345_58_1_n_3214,
       inc_add_1345_58_1_n_3215, inc_add_1345_58_1_n_3220,
       inc_add_1345_58_1_n_3222, inc_add_1345_58_1_n_3229;
  wire inc_add_1345_58_1_n_3230, inc_add_1345_58_1_n_3234,
       inc_add_1345_58_1_n_3236, inc_add_1345_58_1_n_3238,
       inc_add_1345_58_1_n_3242, inc_add_1345_58_1_n_3246,
       inc_add_1345_58_1_n_3248, inc_add_1345_58_1_n_3250;
  wire inc_add_1345_58_1_n_3252, inc_add_1345_58_1_n_3254,
       inc_add_1345_58_1_n_3257, inc_add_1345_58_1_n_3258,
       inc_add_1345_58_1_n_3263, inc_add_1345_58_1_n_3266,
       inc_add_1345_58_1_n_3267, inc_add_1345_58_1_n_3271;
  wire inc_add_1345_58_1_n_3273, inc_add_1345_58_1_n_3279,
       inc_add_1345_58_1_n_3280, inc_add_1345_58_1_n_3283,
       inc_add_1345_58_1_n_3288, inc_add_1345_58_1_n_3293,
       inc_add_1345_58_1_n_3298, inc_add_1345_58_1_n_3301;
  wire inc_add_1345_58_1_n_3304, inc_add_1345_58_1_n_3307,
       inc_add_1345_58_1_n_3310, inc_add_1345_58_1_n_3315,
       inc_add_1345_58_1_n_3320, inc_add_1345_58_1_n_3325,
       inc_add_1345_58_1_n_3330, inc_add_1345_58_1_n_3335;
  wire inc_add_1345_58_1_n_3338, inc_add_1345_58_1_n_3343,
       inc_add_1345_58_1_n_3348, inc_add_1345_58_1_n_3353,
       inc_add_1345_58_1_n_3358, inc_add_1345_58_1_n_3364,
       inc_add_1345_58_1_n_3366, inc_add_1345_58_1_n_3370;
  wire inc_add_1345_58_1_n_3373, inc_add_1345_58_1_n_3378,
       inc_add_1345_58_1_n_3382, inc_add_1345_58_1_n_3387,
       inc_add_1345_58_1_n_3390, inc_add_1345_58_1_n_3399,
       inc_add_1345_58_1_n_3408, inc_add_1345_58_1_n_3414;
  wire inc_add_1345_58_1_n_3422, inc_add_1345_58_1_n_3434,
       inc_add_1345_58_1_n_3455, inc_add_1347_34_2_n_2311,
       inc_add_1347_34_2_n_2316, inc_add_1347_34_2_n_2321,
       inc_add_1347_34_2_n_2326, inc_add_1347_34_2_n_2331;
  wire inc_add_1347_34_2_n_2336, inc_add_1347_34_2_n_2341,
       inc_add_1347_34_2_n_2347, inc_add_1347_34_2_n_2352,
       inc_add_1347_34_2_n_2357, inc_add_1347_34_2_n_2362,
       inc_add_1347_34_2_n_2368, inc_add_1347_34_2_n_2373;
  wire inc_add_1347_34_2_n_2377, inc_add_1347_34_2_n_2381,
       inc_add_1347_34_2_n_2389, inc_add_1347_34_2_n_2391,
       inc_add_1347_34_2_n_2396, inc_add_1347_34_2_n_2400,
       inc_add_1347_34_2_n_2401, inc_add_1347_34_2_n_2409;
  wire inc_add_1347_34_2_n_2411, inc_add_1347_34_2_n_2413,
       inc_add_1347_34_2_n_2417, inc_add_1347_34_2_n_2422,
       inc_add_1347_34_2_n_2426, inc_add_1347_34_2_n_2429,
       inc_add_1347_34_2_n_2431, inc_add_1347_34_2_n_2434;
  wire inc_add_1347_34_2_n_2436, inc_add_1347_34_2_n_2439,
       inc_add_1347_34_2_n_2441, inc_add_1347_34_2_n_2445,
       inc_add_1347_34_2_n_2446, inc_add_1347_34_2_n_2449,
       inc_add_1347_34_2_n_2451, inc_add_1347_34_2_n_2453;
  wire inc_add_1347_34_2_n_2455, inc_add_1347_34_2_n_2457,
       inc_add_1347_34_2_n_2459, inc_add_1347_34_2_n_2461,
       inc_add_1347_34_2_n_2462, inc_add_1347_34_2_n_2464,
       inc_add_1347_34_2_n_2467, inc_add_1347_34_2_n_2472;
  wire inc_add_1347_34_2_n_2482, inc_add_1347_34_2_n_2487,
       inc_add_1347_34_2_n_2492, inc_add_1347_34_2_n_2497,
       inc_add_1347_34_2_n_2502, inc_add_1347_34_2_n_2505,
       inc_add_1347_34_2_n_2510, inc_add_1347_34_2_n_2515;
  wire inc_add_1347_34_2_n_2520, inc_add_1347_34_2_n_2525,
       inc_add_1347_34_2_n_2530, inc_add_1347_34_2_n_2536,
       inc_add_1347_34_2_n_2538, inc_add_1347_34_2_n_2544,
       inc_add_1347_34_2_n_2547, inc_add_1347_34_2_n_2553;
  wire inc_add_1347_34_2_n_2558, inc_add_1347_34_2_n_2561,
       inc_add_1347_34_2_n_2589, inc_add_1347_34_2_n_2595,
       inc_add_1347_34_2_n_2650, inc_add_1347_34_2_n_2652,
       \instruction[5]_40251 , \instruction[7]_39642 ;
  wire \instruction[8]_40127 , \instruction[9]_40095 ,
       \instruction[10]_40063 , \instruction[11]_40312 ,
       \instruction[14]_40189 , \instruction_address[0] , jal_type,
       load_request_BAR;
  wire n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8;
  wire n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16;
  wire n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24;
  wire n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32;
  wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40;
  wire n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_173, n_174, n_175, n_178, n_179;
  wire n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187;
  wire n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195;
  wire n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203;
  wire n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211;
  wire n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219;
  wire n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227;
  wire n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_245, n_246, n_249, n_250, n_251, n_252, n_253;
  wire n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_676, n_677, n_678, n_679, n_680, n_682, n_683;
  wire n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691;
  wire n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_748, n_750, n_751, n_752, n_753, n_754, n_755, n_756;
  wire n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764;
  wire n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772;
  wire n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780;
  wire n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788;
  wire n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796;
  wire n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804;
  wire n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812;
  wire n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820;
  wire n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836;
  wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868;
  wire n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884;
  wire n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892;
  wire n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900;
  wire n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956;
  wire n_957, n_958, n_959, n_960, n_962, n_963, n_964, n_965;
  wire n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973;
  wire n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981;
  wire n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989;
  wire n_990, n_991, n_993, n_994, n_995, n_996, n_997, n_998;
  wire n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006;
  wire n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014;
  wire n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022;
  wire n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030;
  wire n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038;
  wire n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046;
  wire n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054;
  wire n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062;
  wire n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070;
  wire n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078;
  wire n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1088;
  wire n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1105, n_1106;
  wire n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130;
  wire n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146;
  wire n_1147, n_1148, n_1149, n_1150, n_1151, n_1153, n_1154, n_1155;
  wire n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
  wire n_1164, n_1165, n_1166, n_1167, n_1169, n_1170, n_1171, n_1172;
  wire n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180;
  wire n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196;
  wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1205;
  wire n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1214;
  wire n_1216, n_1217, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224;
  wire n_1227, n_1229, n_1230, n_1231, n_1232, n_1233, n_1235, n_1236;
  wire n_1237, n_1239, n_1240, n_1242, n_1243, n_1246, n_1247, n_1249;
  wire n_1250, n_1251, n_1253, n_1254, n_1256, n_1257, n_1258, n_1260;
  wire n_1261, n_1263, n_1264, n_1266, n_1267, n_1268, n_1269, n_1270;
  wire n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278;
  wire n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286;
  wire n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294;
  wire n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302;
  wire n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310;
  wire n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318;
  wire n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326;
  wire n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334;
  wire n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342;
  wire n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350;
  wire n_1351, n_1352, n_1353, n_1354, n_1356, n_1357, n_1358, n_1359;
  wire n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367;
  wire n_1368, n_1369, n_1370, n_1372, n_1373, n_1374, n_1375, n_1376;
  wire n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400;
  wire n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408;
  wire n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416;
  wire n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425;
  wire n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433;
  wire n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441;
  wire n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449;
  wire n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465;
  wire n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473;
  wire n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481;
  wire n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489;
  wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505;
  wire n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513;
  wire n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521;
  wire n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529;
  wire n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537;
  wire n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545;
  wire n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553;
  wire n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561;
  wire n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569;
  wire n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577;
  wire n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585;
  wire n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593;
  wire n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601;
  wire n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609;
  wire n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617;
  wire n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625;
  wire n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633;
  wire n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641;
  wire n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649;
  wire n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657;
  wire n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665;
  wire n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673;
  wire n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681;
  wire n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689;
  wire n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697;
  wire n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705;
  wire n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713;
  wire n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721;
  wire n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729;
  wire n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737;
  wire n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745;
  wire n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753;
  wire n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761;
  wire n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769;
  wire n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777;
  wire n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785;
  wire n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793;
  wire n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801;
  wire n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809;
  wire n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817;
  wire n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825;
  wire n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833;
  wire n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841;
  wire n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849;
  wire n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857;
  wire n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865;
  wire n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873;
  wire n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881;
  wire n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889;
  wire n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897;
  wire n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905;
  wire n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913;
  wire n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921;
  wire n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929;
  wire n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937;
  wire n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945;
  wire n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953;
  wire n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961;
  wire n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969;
  wire n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977;
  wire n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985;
  wire n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993;
  wire n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001;
  wire n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009;
  wire n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017;
  wire n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025;
  wire n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033;
  wire n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041;
  wire n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049;
  wire n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057;
  wire n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065;
  wire n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073;
  wire n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081;
  wire n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089;
  wire n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097;
  wire n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105;
  wire n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113;
  wire n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121;
  wire n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129;
  wire n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137;
  wire n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145;
  wire n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153;
  wire n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161;
  wire n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169;
  wire n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177;
  wire n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185;
  wire n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193;
  wire n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201;
  wire n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209;
  wire n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217;
  wire n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225;
  wire n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233;
  wire n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241;
  wire n_2242, n_2243, n_2244, n_2245, n_2246, n_2248, n_2249, n_2250;
  wire n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258;
  wire n_2259, n_2260, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268;
  wire n_2269, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277;
  wire n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285;
  wire n_2286, n_2287, n_2288, n_2289, n_2290, n_2292, n_2293, n_2294;
  wire n_2295, n_2296, n_2297, n_2298, n_2300, n_2303, n_2304, n_2305;
  wire n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313;
  wire n_2314, n_2316, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323;
  wire n_2324, n_2325, n_2326, n_2328, n_2329, n_2330, n_2331, n_2332;
  wire n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340;
  wire n_2343, n_2345, n_2346, n_2347, n_2348, n_2349, n_2351, n_2352;
  wire n_2353, n_2357, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364;
  wire n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372;
  wire n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380;
  wire n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2388, n_2389;
  wire n_2390, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398;
  wire n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406;
  wire n_2407, n_2408, n_2409, n_2410, n_2411, n_2414, n_2415, n_2416;
  wire n_2417, n_2418, n_2419, n_2420, n_2421, n_2423, n_2424, n_2425;
  wire n_2426, n_2428, n_2429, n_2431, n_2432, n_2433, n_2435, n_2437;
  wire n_2438, n_2439, n_2440, n_2441, n_2442, n_2444, n_2445, n_2446;
  wire n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454;
  wire n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462;
  wire n_2463, n_2464, n_2465, n_2466, n_2467, n_2472, n_2474, n_2475;
  wire n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483;
  wire n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491;
  wire n_2492, n_2493, n_2495, n_2496, n_2497, n_2498, n_2500, n_2501;
  wire n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509;
  wire n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517;
  wire n_2518, n_2520, n_2521, n_2522, n_2523, n_2524, n_2526, n_2527;
  wire n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535;
  wire n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543;
  wire n_2544, n_2545, n_2546, n_2548, n_2549, n_2550, n_2551, n_2552;
  wire n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560;
  wire n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568;
  wire n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2576, n_2577;
  wire n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585;
  wire n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593;
  wire n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602;
  wire n_2603, n_2604, n_2606, n_2609, n_2611, n_2613, n_2614, n_2615;
  wire n_2619, n_2620, n_2621, n_2622, n_2623, n_2625, n_2626, n_2627;
  wire n_2628, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636;
  wire n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2644, n_2645;
  wire n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2653, n_2654;
  wire n_2655, n_2656, n_2658, n_2659, n_2660, n_2661, n_2662, n_2664;
  wire n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2676;
  wire n_2678, n_2680, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687;
  wire n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695;
  wire n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703;
  wire n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711;
  wire n_2712, n_2713, n_2714, n_2715, n_2718, n_2719, n_2720, n_2721;
  wire n_2722, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2731;
  wire n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739;
  wire n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748;
  wire n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756;
  wire n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764;
  wire n_2765, n_2766, n_2767, n_2768, n_2771, n_2772, n_2773, n_2774;
  wire n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782;
  wire n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791;
  wire n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799;
  wire n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2807, n_2808;
  wire n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816;
  wire n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824;
  wire n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832;
  wire n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840;
  wire n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848;
  wire n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856;
  wire n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864;
  wire n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872;
  wire n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880;
  wire n_2881, n_2882, n_2883, n_2884, n_2885, n_2887, n_2888, n_2889;
  wire n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897;
  wire n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905;
  wire n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913;
  wire n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921;
  wire n_2922, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, n_2930;
  wire n_2931, n_2932, n_2933, n_2934, n_2936, n_2937, n_2938, n_2939;
  wire n_2940, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948;
  wire n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956;
  wire n_2957, n_2958, n_2959, n_2960, n_2962, n_2963, n_2964, n_2965;
  wire n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973;
  wire n_2975, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983;
  wire n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991;
  wire n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999;
  wire n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007;
  wire n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015;
  wire n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023;
  wire n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031;
  wire n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039;
  wire n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047;
  wire n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055;
  wire n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063;
  wire n_3064, n_3065, n_3066, n_3069, n_3071, n_3073, n_3074, n_3075;
  wire n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083;
  wire n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091;
  wire n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099;
  wire n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107;
  wire n_3108, n_3109, n_3110, n_3112, n_3113, n_3114, n_3115, n_3117;
  wire n_3118, n_3119, n_3123, n_3126, n_3127, n_3129, n_3130, n_3131;
  wire n_3132, n_3133, n_3134, n_3135, n_3137, n_3138, n_3140, n_3141;
  wire n_3142, n_3145, n_3147, n_3149, n_3150, n_3151, n_3152, n_3153;
  wire n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161;
  wire n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169;
  wire n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177;
  wire n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3186;
  wire n_3187, n_3188, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195;
  wire n_3196, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204;
  wire n_3205, n_3206, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213;
  wire n_3214, n_3215, n_3216, n_3217, n_3218, n_3220, n_3221, n_3222;
  wire n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3230, n_3231;
  wire n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239;
  wire n_3240, n_3241, n_3242, n_3243, n_3245, n_3246, n_3247, n_3248;
  wire n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3257, n_3259;
  wire n_3260, n_3261, n_3262, n_3263, n_3264, n_3266, n_3267, n_3268;
  wire n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277;
  wire n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287;
  wire n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295;
  wire n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303;
  wire n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311;
  wire n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3320;
  wire n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328;
  wire n_3329, n_3330, n_3331, n_3335, n_3336, n_3337, n_3338, n_3340;
  wire n_3341, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350;
  wire n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358;
  wire n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366;
  wire n_3367, n_3373, n_3374, n_3375, n_3376, n_3378, n_3379, n_3380;
  wire n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388;
  wire n_3389, n_3390, n_3391, n_3392, n_3393, n_3395, n_3396, n_3397;
  wire n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405;
  wire n_3406, n_3407, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414;
  wire n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422;
  wire n_3423, n_3424, n_3426, n_3427, n_3428, n_3429, n_3431, n_3432;
  wire n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440;
  wire n_3441, n_3442, n_3444, n_3445, n_3449, n_3450, n_3451, n_3452;
  wire n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460;
  wire n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3468, n_3469;
  wire n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477;
  wire n_3478, n_3479, n_3480, n_3482, n_3483, n_3484, n_3485, n_3486;
  wire n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494;
  wire n_3495, n_3496, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503;
  wire n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511;
  wire n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519;
  wire n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527;
  wire n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535;
  wire n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543;
  wire n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551;
  wire n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559;
  wire n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567;
  wire n_3570, n_3572, n_3573, n_3574, n_3576, n_3578, n_3579, n_3580;
  wire n_3581, n_3582, n_3583, n_3584, n_3587, n_3588, n_3589, n_3590;
  wire n_3591, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599;
  wire n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607;
  wire n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615;
  wire n_3616, n_3617, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625;
  wire n_3626, n_3628, n_3629, n_3631, n_3632, n_3633, n_3634, n_3635;
  wire n_3636, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3646;
  wire n_3647, n_3648, n_3651, n_3652, n_3653, n_3655, n_3657, n_3658;
  wire n_3660, n_3661, n_3662, n_3663, n_3664, n_3666, n_3667, n_3669;
  wire n_3670, n_3671, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680;
  wire n_3681, n_3682, n_3683, n_3685, n_3686, n_3687, n_3688, n_3689;
  wire n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3697, n_3698;
  wire n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706;
  wire n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714;
  wire n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722;
  wire n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730;
  wire n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738;
  wire n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746;
  wire n_3747, n_3748, n_3750, n_3752, n_3753, n_3755, n_3756, n_3757;
  wire n_3758, n_3759, n_3760, n_3761, n_3763, n_3764, n_3766, n_3767;
  wire n_3768, n_3770, n_3773, n_3777, n_3778, n_3779, n_3780, n_3781;
  wire n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793;
  wire n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801;
  wire n_3802, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810;
  wire n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818;
  wire n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826;
  wire n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834;
  wire n_3835, n_3836, n_3838, n_3839, n_3841, n_3842, n_3845, n_3846;
  wire n_3848, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856;
  wire n_3857, n_3858, n_3859, n_3860, n_3862, n_3863, n_3864, n_3866;
  wire n_3869_BAR, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876,
       n_3877;
  wire n_3880, n_3881, n_3882, n_3883, n_3884, n_3886, n_3887, n_3888;
  wire n_3891, n_3892, n_3893, n_3894, n_3897, n_3898, n_3899, n_3900;
  wire n_3902, n_3905, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912;
  wire n_3913, n_3915, n_3916, n_3917, n_3918, n_3920, n_3921, n_3922;
  wire n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930;
  wire n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938;
  wire n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946;
  wire n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953, n_3954;
  wire n_3955, n_3956, n_3957, n_3958, n_3961, n_3962, n_3963, n_3964;
  wire n_3965, n_3966, n_3967, n_3968, n_3969, n_3971, n_3972, n_3973;
  wire n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982, n_3983;
  wire n_3984, n_3986, n_3987, n_3988, n_3989, n_3990, n_3992, n_3993;
  wire n_3994, n_3995, n_3996, n_3999, n_4000, n_4001, n_4002, n_4007;
  wire n_4008, n_4009, n_4010, n_4011, n_4013, n_4014, n_4015, n_4016;
  wire n_4017, n_4018, n_4019, n_4021, n_4022, n_4023, n_4024, n_4025;
  wire n_4026, n_4027, n_4028, n_4030, n_4031, n_4032, n_4033, n_4035;
  wire n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, n_4043;
  wire n_4044, n_4045, n_4046, n_4048, n_4049, n_4050, n_4051, n_4052;
  wire n_4053, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, n_4061;
  wire n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069;
  wire n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077;
  wire n_4078, n_4079, n_4080, n_4082, n_4083, n_4084, n_4085, n_4087;
  wire n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095;
  wire n_4096, n_4097, n_4100, n_4101, n_4102, n_4103, n_4104, n_4107;
  wire n_4108, n_4109, n_4111, n_4112, n_4114, n_4115, n_4116, n_4118;
  wire n_4119, n_4121, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128;
  wire n_4129, n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4137;
  wire n_4138, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145, n_4146;
  wire n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153, n_4154;
  wire n_4155, n_4156, n_4159, n_4161, n_4162, n_4164, n_4165, n_4166;
  wire n_4167, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174, n_4175;
  wire n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182, n_4185;
  wire n_4186, n_4187, n_4188, n_4189, n_4190, n_4192, n_4193, n_4194;
  wire n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201, n_4202;
  wire n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4210, n_4212;
  wire n_4213, n_4214, n_4215, n_4221, n_4223, n_4224, n_4225, n_4226;
  wire n_4227, n_4228, n_4229, n_4230, n_4231, n_4232, n_4234, n_4235;
  wire n_4236, n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243;
  wire n_4244, n_4245, n_4246, n_4247, n_4249, n_4250, n_4251, n_4252;
  wire n_4253, n_4254, n_4255, n_4256, n_4262, n_4263, n_4264, n_4267;
  wire n_4268, n_4270, n_4272, n_4273, n_4274, n_4277, n_4278, n_4279;
  wire n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291;
  wire n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, n_4299;
  wire n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308;
  wire n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317;
  wire n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325;
  wire n_4326, n_4328, n_4329, n_4330, n_4331, n_4332, n_4333, n_4334;
  wire n_4335, n_4336, n_4337, n_4338, n_4339, n_4340, n_4341, n_4342;
  wire n_4343, n_4344, n_4345, n_4346, n_4347, n_4348, n_4349, n_4350;
  wire n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357, n_4358;
  wire n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, n_4366, n_4367;
  wire n_4368, n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375;
  wire n_4376, n_4377, n_4378, n_4379, n_4380, n_4381, n_4382, n_4383;
  wire n_4384, n_4385, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391;
  wire n_4392, n_4393, n_4394, n_4395, n_4396, n_4397, n_4398, n_4399;
  wire n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407;
  wire n_4408, n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415;
  wire n_4416, n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423;
  wire n_4424, n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431;
  wire n_4432, n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439;
  wire n_4440, n_4441, n_4442, n_4443, n_4444, n_4445, n_4446, n_4447;
  wire n_4448, n_4449, n_4450, n_4451, n_4452, n_4453, n_4454, n_4455;
  wire n_4456, n_4457, n_4458, n_4459, n_4460, n_4462, n_4463, n_4464;
  wire n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472;
  wire n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4480, n_4481;
  wire n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488, n_4489;
  wire n_4490, n_4491, n_4492, n_4494, n_4497, n_4498, n_4499, n_4500;
  wire n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509;
  wire n_4510, n_4511, n_4517, n_4522, n_4523, n_4525, n_4526, n_4527;
  wire n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534, n_4535;
  wire n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4543;
  wire n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551;
  wire n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559;
  wire n_4560, n_4561, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567;
  wire n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575;
  wire n_4576, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584;
  wire n_4585, n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592;
  wire n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600;
  wire n_4601, n_4608, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616;
  wire n_4617, n_4620, n_4622, n_4627, n_4628, n_4629, n_4630, n_4631;
  wire n_4632, n_4633, n_4634, n_4636, n_4637, n_4638, n_4639, n_4640;
  wire n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4648, n_4649;
  wire n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658;
  wire n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4666, n_4667;
  wire n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4675;
  wire n_4676, n_4677, n_4678, n_4679, n_4680, n_4682, n_4683, n_4684;
  wire n_4685, n_4686, n_4687, n_4688, n_4689, n_4690, n_4691, n_4692;
  wire n_4693, n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700;
  wire n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, n_4708;
  wire n_4710, n_4711, n_4712, n_4713, n_4714, n_4715, n_4716, n_4717;
  wire n_4718, n_4719, n_4720, n_4723, n_4724, n_4725, n_4726, n_4727;
  wire n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734, n_4735;
  wire n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742, n_4743;
  wire n_4744, n_4745, n_4747, n_4748, n_4750, n_4751, n_4752, n_4753;
  wire n_4755, n_4756, n_4759, n_4761, n_4762, n_4763, n_4764, n_4765;
  wire n_4766, n_4768, n_4769, n_4773, n_4774, n_4775, n_4776, n_4777;
  wire n_4778, n_4781, n_4782, n_4783, n_4784, n_4785, n_4786, n_4787;
  wire n_4788, n_4789, n_4790, n_4791, n_4792, n_4793, n_4794, n_4795;
  wire n_4796, n_4797, n_4798, n_4800, n_4803, n_4804, n_4805, n_4807;
  wire n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815;
  wire n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822, n_4823;
  wire n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831;
  wire n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839;
  wire n_4840, n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847;
  wire n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855;
  wire n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863;
  wire n_4865, n_4866, n_4868, n_4869, n_4870, n_4871, n_4873, n_4874;
  wire n_4876, n_4877, n_4878, n_4879, n_4880, n_4881, n_4882, n_4883;
  wire n_4884, n_4885, n_4886, n_4887, n_4888, n_4889, n_4891, n_4892;
  wire n_4893, n_4894, n_4895, n_4896, n_4897, n_4898, n_4899, n_4900;
  wire n_4901, n_4902, n_4903, n_4904, n_4905, n_4906, n_4907, n_4908;
  wire n_4909, n_4910, n_4911, n_4912, n_4913, n_4914, n_4915, n_4916;
  wire n_4917, n_4918, n_4919, n_4920, n_4921, n_4922, n_4923, n_4924;
  wire n_4925, n_4926, n_4927, n_4928, n_4929, n_4930, n_4931, n_4932;
  wire n_4933, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944;
  wire n_4945, n_4946, n_4947, n_4948, n_4949, n_4952, n_4953, n_4954;
  wire n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4962;
  wire n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970;
  wire n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978;
  wire n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986;
  wire n_4987, n_4988, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994;
  wire n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003;
  wire n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011;
  wire n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019;
  wire n_5020, n_5021, n_5024, n_5025, n_5026, n_5027, n_5028, n_5029;
  wire n_5030, n_5031, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039;
  wire n_5040, n_5041, n_5042, n_5043, n_5044, n_5045, n_5046, n_5047;
  wire n_5048, n_5050, n_5051, n_5053, n_5054, n_5055, n_5058, n_5060;
  wire n_5061, n_5062, n_5066, n_5067, n_5068, n_5070, n_5071, n_5072;
  wire n_5073, n_5075, n_5076, n_5078, n_5079, n_5080, n_5082, n_5083;
  wire n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091;
  wire n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5099, n_5100;
  wire n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108;
  wire n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116;
  wire n_5121, n_5122, n_5123, n_5124, n_5125, n_5126, n_5127, n_5128;
  wire n_5129, n_5130, n_5131, n_5132, n_5133, n_5134, n_5135, n_5136;
  wire n_5137, n_5140, n_5141, n_5143, n_5145, n_5146, n_5147, n_5148;
  wire n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155, n_5156;
  wire n_5157, n_5159, n_5160, n_5161, n_5162, n_5163, n_5164, n_5165;
  wire n_5166, n_5167, n_5168, n_5169, n_5170, n_5171, n_5172, n_5173;
  wire n_5174, n_5175, n_5176, n_5177, n_5178, n_5179, n_5180, n_5181;
  wire n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5190, n_5191;
  wire n_5192, n_5193, n_5194, n_5195, n_5196, n_5197, n_5198, n_5199;
  wire n_5200, n_5201, n_5202, n_5204, n_5205, n_5206, n_5207, n_5208;
  wire n_5209, n_5210, n_5211, n_5213, n_5214, n_5215, n_5216, n_5217;
  wire n_5220, n_5221, n_5222, n_5223, n_5224, n_5225, n_5227, n_5228;
  wire n_5229, n_5230, n_5241, n_5242, n_5243, n_5244, n_5247, n_5248;
  wire n_5249, n_5250, n_5251, n_5252, n_5254, n_5255, n_5256, n_5257;
  wire n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5267;
  wire n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275;
  wire n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283;
  wire n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5292, n_5294;
  wire n_5295, n_5296, n_5297, n_5298, n_5299, n_5300, n_5301, n_5302;
  wire n_5303, n_5304, n_5305, n_5306, n_5307, n_5308, n_5309, n_5312;
  wire n_5313, n_5314, n_5315, n_5320, n_5321, n_5324, n_5325, n_5326;
  wire n_5328, n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335;
  wire n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343;
  wire n_5345, n_5346, n_5347, n_5349, n_5350, n_5351, n_5352, n_5353;
  wire n_5354, n_5357, n_5358, n_5359, n_5362, n_5366, n_5367, n_5368;
  wire n_5371, n_5372, n_5373, n_5374, n_5375, n_5376, n_5377, n_5378;
  wire n_5379, n_5380, n_5381, n_5382, n_5383, n_5387, n_5388, n_5389;
  wire n_5390, n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397;
  wire n_5398, n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405;
  wire n_5406, n_5407, n_5408, n_5409, n_5410, n_5412, n_5413, n_5416;
  wire n_5417, n_5418, n_5419, n_5421, n_5422, n_5423, n_5424, n_5426;
  wire n_5427, n_5430, n_5431, n_5432, n_5434, n_5435, n_5438, n_5440;
  wire n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5449, n_5450;
  wire n_5451, n_5452, n_5453, n_5454, n_5456, n_5458, n_5459, n_5460;
  wire n_5461, n_5462, n_5463, n_5464, n_5465, n_5466, n_5468, n_5469;
  wire n_5472, n_5474, n_5475, n_5476, n_5477, n_5478, n_5480, n_5481;
  wire n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488, n_5489;
  wire n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5500, n_5501;
  wire n_5502, n_5503, n_5504, n_5505, n_5507, n_5508, n_5509, n_5510;
  wire n_5511, n_5512, n_5513, n_5514, n_5516, n_5518, n_5519, n_5520;
  wire n_5521, n_5522, n_5523, n_5524, n_5526, n_5527, n_5528, n_5529;
  wire n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536, n_5538;
  wire n_5539, n_5540, n_5541, n_5542, n_5544, n_5545, n_5546, n_5547;
  wire n_5548, n_5549, n_5550, n_5551, n_5552, n_5553, n_5554, n_5555;
  wire n_5556, n_5557, n_5558, n_5559, n_5560, n_5561, n_5562, n_5563;
  wire n_5564, n_5565, n_5566, n_5567, n_5569, n_5570, n_5571, n_5572;
  wire n_5573, n_5574, n_5575, n_5576, n_5578, n_5579, n_5581, n_5582;
  wire n_5583, n_5584, n_5585, n_5591, n_5593, n_5594, n_5595, n_5598;
  wire n_5599, n_5600, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607;
  wire n_5608, n_5609, n_5610, n_5611, n_5612, n_5613, n_5614, n_5615;
  wire n_5616, n_5617, n_5618, n_5619, n_5620, n_5623, n_5624, n_5626;
  wire n_5627, n_5629, n_5630, n_5632, n_5633, n_5634, n_5635, n_5637;
  wire n_5638, n_5639, n_5640, n_5641, n_5642, n_5644, n_5645, n_5646;
  wire n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653, n_5655;
  wire n_5656, n_5657, n_5658, n_5659, n_5660, n_5661, n_5662, n_5663;
  wire n_5665, n_5666, n_5667, n_5668, n_5669, n_5670, n_5671, n_5672;
  wire n_5674, n_5675, n_5677, n_5678, n_5680, n_5681, n_5683, n_5684;
  wire n_5686, n_5688, n_5689, n_5690, n_5692, n_5693, n_5694, n_5695;
  wire n_5696, n_5697, n_5698, n_5702, n_5704, n_5705, n_5706, n_5707;
  wire n_5708, n_5709, n_5710, n_5711, n_5713, n_5714, n_5715, n_5716;
  wire n_5717, n_5718, n_5719, n_5720, n_5721, n_5723, n_5724, n_5725;
  wire n_5726, n_5727, n_5728, n_5729, n_5730, n_5731, n_5733, n_5734;
  wire n_5735, n_5736, n_5737, n_5738, n_5739, n_5741, n_5744, n_5745;
  wire n_5747, n_5748, n_5754, n_5756, n_5761, n_5764, n_5765, n_5766;
  wire n_5767, n_5768, n_5770, n_5771, n_5772, n_5773, n_5774, n_5776;
  wire n_5777, n_5781, n_5782, n_5784, n_5785, n_5786, n_5787, n_5788;
  wire n_5789, n_5790, n_5791, n_5792, n_5793, n_5795, n_5796, n_5797;
  wire n_5798, n_5799, n_5801, n_5803, n_5804, n_5805, n_5806, n_5807;
  wire n_5808, n_5815, n_5816, n_5819, n_5820, n_5821, n_5822, n_5823;
  wire n_5824, n_5825, n_5826, n_5828, n_5831, n_5837, n_5840, n_5841;
  wire n_5842, n_5843, n_5845, n_5847, n_5848, n_5851, n_5855, n_5856;
  wire n_5857, n_5858, n_5862, n_5863, n_5868, n_5869, n_5870, n_5871;
  wire n_5873, n_5875, n_5877, n_5878, n_5879, n_5880, n_5881, n_5884;
  wire n_5885, n_5886, n_5887, n_5892, n_5893, n_5903, n_5904, n_5906;
  wire n_5907, n_5911, n_5919, n_5924, n_5927, n_5930, n_5932, n_5933;
  wire n_5935, n_5936, n_5938, n_5941, n_5942, n_5945, n_5947, n_5950;
  wire n_5951, n_5955, n_5956, n_5957, n_5958, n_5959, n_5961, n_5962;
  wire n_5963, n_5964, n_5965, n_5972, n_5973, n_5975, n_5976, n_5978;
  wire n_5979, n_5980, n_5984, n_5986, n_5989, n_5990, n_5991, n_5992;
  wire n_5994, n_5995, n_5996, n_5998, n_6000, n_6003, n_6006, n_6007;
  wire n_6008, n_6009, n_6011, n_6012, n_6013, n_6015, n_6017, n_6022;
  wire n_6023, n_6024, n_6025, n_6026, n_6027, n_6028, n_6033, n_6034;
  wire n_6035, n_6036, n_6037, n_6038, n_6039, n_6040, n_6041, n_6042;
  wire n_6043, n_6044, n_6045, n_6046, n_6047, n_6048, n_6049, n_6050;
  wire n_6052, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6060;
  wire n_6061, n_6062, n_6064, n_6065, n_6066, n_6067, n_6068, n_6070;
  wire n_6071, n_6072, n_6073, n_6074, n_6075, n_6076, n_6077, n_6078;
  wire n_6079, n_6080, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087;
  wire n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095;
  wire n_6096, n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103;
  wire n_6104, n_6105, n_6106, n_6107, n_6108, n_6109, n_6110, n_6111;
  wire n_6112, n_6113, n_6114, n_6121, n_6123, n_6126, n_6127, n_6132;
  wire n_6134, n_6135, n_6136, n_6137, n_6139, n_6141, n_6143, n_6145;
  wire n_6149, n_6153, n_6155, n_6159, n_6161, n_6165, n_6167, n_6170;
  wire n_6178, n_6181, n_6183, n_6195, n_6232, n_6233, n_6234, n_6235;
  wire n_6236, n_6237, n_6238, n_6256, n_6257, n_6258, n_6259, n_6260;
  wire n_6261, n_6262, n_6263, n_6264, n_6265, n_6266, n_6267, n_6268;
  wire n_6269, n_6270, n_6271, n_6272, n_6273, n_6274, n_6275, n_6276;
  wire n_6277, n_6278, n_6279, n_6280, n_6281, n_6282, n_6283, n_6284;
  wire n_6285, n_6286, n_6287, n_6288, n_6289, n_6290, n_6291, n_6292;
  wire n_6293, n_6294, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300;
  wire n_6301, n_6302, n_6303, n_6304, n_6305, n_6306, n_6307, n_6308;
  wire n_6309, n_6310, n_6311, n_6312, n_6313, n_6314, n_6315, n_6316;
  wire n_6317, n_6318, n_6319, n_6320, n_6321, n_6322, n_6323, n_6324;
  wire n_6325, n_6326, n_6327, n_6328, n_6329, n_6330, n_6331, n_6332;
  wire n_6333, n_6334, n_6335, n_6336, n_6337, n_6338, n_6339, n_6340;
  wire n_6341, n_6342, n_6343, n_6344, n_6345, n_6346, n_6347, n_6348;
  wire n_6349, n_6350, n_6351, n_6352, n_6353, n_6354, n_6355, n_6356;
  wire n_6357, n_6358, n_6359, n_6360, n_6361, n_6362, n_6363, n_6364;
  wire n_6365, n_6366, n_6367, n_6368, n_6369, n_6370, n_6371, n_6372;
  wire n_6373, n_6374, n_6375, n_6376, n_6377, n_6378, n_6379, n_6380;
  wire n_6381, n_6382, n_6383, n_6384, n_6385, n_6386, n_6387, n_6388;
  wire n_6389, n_6390, n_6391, n_6392, n_6393, n_6394, n_6395, n_6396;
  wire n_6397, n_6398, n_6399, n_6400, n_6401, n_6402, n_6403, n_6404;
  wire n_6405, n_6406, n_6407, n_6408, n_6409, n_6410, n_6411, n_6412;
  wire n_6413, n_6414, n_6415, n_6416, n_6417, n_6418, n_6419, n_6420;
  wire n_6421, n_6422, n_6423, n_6424, n_6425, n_6426, n_6427, n_6428;
  wire n_6429, n_6430, n_6431, n_6432, n_6433, n_6434, n_6435, n_6436;
  wire n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443, n_6444;
  wire n_6445, n_6446, n_6447, n_6448, n_6449, n_6450, n_6451, n_6452;
  wire n_6453, n_6454, n_6455, n_6456, n_6457, n_6458, n_6459, n_6460;
  wire n_6461, n_6462, n_6463, n_6464, n_6465, n_6466, n_6467, n_6468;
  wire n_6469, n_6470, n_6471, n_6472, n_6473, n_6474, n_6475, n_6476;
  wire n_6477, n_6478, n_6479, n_6480, n_6481, n_6482, n_6483, n_6484;
  wire n_6485, n_6486, n_6487, n_6488, n_6489, n_6490, n_6491, n_6492;
  wire n_6493, n_6494, n_6495, n_6496, n_6497, n_6498, n_6499, n_6500;
  wire n_6501, n_6502, n_6503, n_6504, n_6505, n_6506, n_6507, n_6508;
  wire n_6509, n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6516;
  wire n_6517, n_6518, n_6519, n_6520, n_6521, n_6522, n_6523, n_6524;
  wire n_6525, n_6526, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532;
  wire n_6533, n_6534, n_6535, n_6536, n_6537, n_6538, n_6539, n_6540;
  wire n_6541, n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548;
  wire n_6549, n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556;
  wire n_6557, n_6558, n_6559, n_6560, n_6561, n_6562, n_6563, n_6564;
  wire n_6565, n_6566, n_6567, n_6568, n_6569, n_6570, n_6571, n_6572;
  wire n_6573, n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, n_6580;
  wire n_6581, n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6588;
  wire n_6589, n_6590, n_6591, n_6592, n_6593, n_6594, n_6595, n_6596;
  wire n_6597, n_6598, n_6599, n_6600, n_6601, n_6602, n_6603, n_6604;
  wire n_6605, n_6606, n_6607, n_6608, n_6609, n_6610, n_6611, n_6612;
  wire n_6613, n_6614, n_6615, n_6616, n_6617, n_6618, n_6619, n_6620;
  wire n_6621, n_6622, n_6623, n_6624, n_6625, n_6626, n_6627, n_6628;
  wire n_6629, n_6630, n_6631, n_6632, n_6633, n_6634, n_6635, n_6636;
  wire n_6637, n_6638, n_6639, n_6640, n_6641, n_6642, n_6643, n_6644;
  wire n_6645, n_6646, n_6647, n_6648, n_6649, n_6650, n_6651, n_6652;
  wire n_6653, n_6654, n_6655, n_6656, n_6657, n_6658, n_6659, n_6660;
  wire n_6661, n_6662, n_6663, n_6664, n_6665, n_6666, n_6667, n_6668;
  wire n_6669, n_6670, n_6671, n_6672, n_6673, n_6674, n_6675, n_6676;
  wire n_6677, n_6678, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684;
  wire n_6685, n_6686, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692;
  wire n_6693, n_6694, n_6695, n_6696, n_6697, n_6698, n_6699, n_6700;
  wire n_6701, n_6702, n_6703, n_6704, n_6705, n_6706, n_6707, n_6708;
  wire n_6709, n_6710, n_6711, n_6712, n_6713, n_6714, n_6715, n_6716;
  wire n_6717, n_6718, n_6719, n_6720, n_6721, n_6722, n_6723, n_6724;
  wire n_6725, n_6726, n_6727, n_6728, n_6729, n_6730, n_6731, n_6732;
  wire n_6733, n_6734, n_6735, n_6736, n_6737, n_6738, n_6739, n_6740;
  wire n_6741, n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748;
  wire n_6749, n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756;
  wire n_6757, n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764;
  wire n_6765, n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772;
  wire n_6773, n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780;
  wire n_6781, n_6782, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788;
  wire n_6789, n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796;
  wire n_6797, n_6798, n_6799, n_6800, n_6801, n_6802, n_6803, n_6804;
  wire n_6805, n_6806, n_6807, n_6808, n_6809, n_6810, n_6811, n_6812;
  wire n_6813, n_6814, n_6815, n_6816, n_6817, n_6818, n_6819, n_6820;
  wire n_6821, n_6822, n_6823, n_6824, n_6825, n_6826, n_6827, n_6828;
  wire n_6829, n_6830, n_6831, n_6832, n_6833, n_6834, n_6835, n_6836;
  wire n_6837, n_6838, n_6839, n_6840, n_6841, n_6842, n_6843, n_6844;
  wire n_6845, n_6846, n_6847, n_6848, n_6849, n_6850, n_6851, n_6852;
  wire n_6853, n_6854, n_6855, n_6856, n_6857, n_6858, n_6859, n_6860;
  wire n_6861, n_6862, n_6863, n_6864, n_6865, n_6866, n_6867, n_6868;
  wire n_6869, n_6870, n_6871, n_6872, n_6873, n_6874, n_6875, n_6876;
  wire n_6877, n_6878, n_6879, n_6880, n_6881, n_6882, n_6883, n_6884;
  wire n_6885, n_6886, n_6887, n_6888, n_6889, n_6890, n_6891, n_6892;
  wire n_6893, n_6894, n_6895, n_6896, n_6897, n_6898, n_6899, n_6900;
  wire n_6901, n_6902, n_6903, n_6904, n_6905, n_6906, n_6907, n_6908;
  wire n_6909, n_6910, n_6911, n_6912, n_6913, n_6914, n_6915, n_6916;
  wire n_6917, n_6918, n_6919, n_6920, n_6921, n_6922, n_6923, n_6924;
  wire n_6925, n_6926, n_6927, n_6928, n_6929, n_6930, n_6931, n_6932;
  wire n_6933, n_6934, n_6935, n_6936, n_6937, n_6938, n_6939, n_6940;
  wire n_6941, n_6942, n_6943, n_6944, n_6945, n_6946, n_6947, n_6948;
  wire n_6949, n_6950, n_6951, n_6952, n_6953, n_6954, n_6955, n_6956;
  wire n_6957, n_6958, n_6959, n_6960, n_6961, n_6962, n_6963, n_6964;
  wire n_6965, n_6966, n_6967, n_6968, n_6969, n_6970, n_6971, n_6972;
  wire n_6973, n_6974, n_6975, n_6976, n_6977, n_6978, n_6979, n_6980;
  wire n_6981, n_6982, n_6983, n_6984, n_6985, n_6986, n_6987, n_6988;
  wire n_6989, n_6990, n_6991, n_6992, n_6993, n_6994, n_6995, n_6996;
  wire n_6997, n_6998, n_6999, n_7000, n_7001, n_7002, n_7003, n_7004;
  wire n_7005, n_7006, n_7007, n_7008, n_7009, n_7010, n_7011, n_7012;
  wire n_7013, n_7014, n_7015, n_7016, n_7017, n_7018, n_7019, n_7020;
  wire n_7021, n_7022, n_7023, n_7024, n_7025, n_7026, n_7027, n_7028;
  wire n_7029, n_7030, n_7031, n_7032, n_7033, n_7034, n_7035, n_7036;
  wire n_7037, n_7038, n_7039, n_7040, n_7041, n_7042, n_7043, n_7044;
  wire n_7045, n_7046, n_7047, n_7048, n_7049, n_7050, n_7051, n_7052;
  wire n_7053, n_7054, n_7055, n_7056, n_7057, n_7058, n_7059, n_7060;
  wire n_7061, n_7062, n_7063, n_7064, n_7065, n_7066, n_7067, n_7068;
  wire n_7069, n_7070, n_7071, n_7072, n_7073, n_7074, n_7075, n_7076;
  wire n_7077, n_7078, n_7079, n_7080, n_7081, n_7082, n_7083, n_7084;
  wire n_7085, n_7086, n_7087, n_7088, n_7089, n_7090, n_7091, n_7092;
  wire n_7093, n_7094, n_7095, n_7096, n_7097, n_7098, n_7099, n_7100;
  wire n_7101, n_7102, n_7103, n_7104, n_7105, n_7106, n_7107, n_7108;
  wire n_7109, n_7110, n_7111, n_7112, n_7113, n_7114, n_7115, n_7116;
  wire n_7117, n_7118, n_7119, n_7120, n_7121, n_7122, n_7123, n_7124;
  wire n_7125, n_7126, n_7127, n_7128, n_7129, n_7130, n_7131, n_7132;
  wire n_7133, n_7134, n_7135, n_7136, n_7137, n_7138, n_7139, n_7140;
  wire n_7141, n_7142, n_7143, n_7144, n_7145, n_7146, n_7147, n_7148;
  wire n_7149, n_7150, n_7151, n_7152, n_7153, n_7154, n_7155, n_7156;
  wire n_7157, n_7158, n_7159, n_7160, n_7161, n_7162, n_7163, n_7164;
  wire n_7165, n_7166, n_7167, n_7168, n_7169, n_7170, n_7171, n_7172;
  wire n_7173, n_7174, n_7175, n_7176, n_7177, n_7178, n_7179, n_7180;
  wire n_7181, n_7182, n_7183, n_7184, n_7185, n_7186, n_7187, n_7188;
  wire n_7189, n_7190, n_7191, n_7192, n_7193, n_7194, n_7195, n_7196;
  wire n_7197, n_7198, n_7199, n_7200, n_7201, n_7202, n_7203, n_7204;
  wire n_7205, n_7206, n_7207, n_7208, n_7209, n_7210, n_7211, n_7212;
  wire n_7213, n_7214, n_7215, n_7216, n_7217, n_7218, n_7219, n_7220;
  wire n_7221, n_7222, n_7223, n_7224, n_7225, n_7226, n_7227, n_7228;
  wire n_7229, n_7230, n_7231, n_7232, n_7233, n_7234, n_7235, n_7236;
  wire n_7237, n_7238, n_7239, n_7240, n_7241, n_7242, n_7243, n_7244;
  wire n_7245, n_7246, n_7247, n_7248, n_7249, n_7250, n_7251, n_7252;
  wire n_7253, n_7254, n_7255, n_7256, n_7257, n_7258, n_7259, n_7260;
  wire n_7261, n_7262, n_7263, n_7264, n_7265, n_7266, n_7267, n_7268;
  wire n_7269, n_7270, n_7271, n_7272, n_7273, n_7274, n_7275, n_7276;
  wire n_7277, n_7278, n_7279, n_7280, n_7282, n_7302, n_7303, n_7304;
  wire n_7305, n_7370, n_7371, n_7376, n_7377, n_7378, n_7379, n_7380;
  wire n_7381, n_7383, n_7384, n_7385, n_7386, n_7387, n_7388, n_7389;
  wire n_7391, n_7392, n_7393, n_7394, n_7395, n_7397, n_7398, n_7399;
  wire n_7400, n_7401, n_7404, n_7406, n_7407, n_7408, n_7409, n_7410;
  wire n_7412, n_7413, n_7414, n_7415, n_7416, n_7417, n_7418, n_7419;
  wire n_7420, n_7421, n_7422, n_7423, n_7424, n_7425, n_7426, n_7427;
  wire n_7428, n_7429, n_7431, n_7433, n_7435, n_7437, n_7438, n_7439;
  wire n_7440, n_7441, n_7442, n_7443, n_7444, n_7445, n_7446, n_7447;
  wire n_7448, n_7449, n_7450, n_7451, n_7452, n_7453, n_7454, n_7455;
  wire n_7456, n_7457, n_7458, n_7459, n_7460, n_7461, n_7462, n_7463;
  wire n_7464, n_7465, n_7467, n_7468, n_7469, n_7470, n_7471, n_7472;
  wire n_7474, n_7475, n_7476, n_7477, n_7478, n_7479, n_7480, n_7481;
  wire n_7482, n_7483, n_7484, n_7485, n_7486, n_7487, n_7488, n_7489;
  wire n_7490, n_7491, n_7492, n_7493, n_7494, n_7495, n_7496, n_7497;
  wire n_7498, n_7499, n_7500, n_7501, n_7502, n_7503, n_7504, n_7505;
  wire n_7506, n_7507, n_7508, n_7509, n_7510, n_7511, n_7512, n_7513;
  wire n_7514, n_7515, n_7516, n_7517, n_7518, n_7519, n_7520, n_7521;
  wire n_7522, n_7523, n_7524, n_7525, n_7526, n_7527, n_7528, n_7529;
  wire n_7530, n_7531, n_7532, n_7533, n_7534, n_7535, n_7536, n_7537;
  wire n_7538, n_7539, n_7540, n_7541, n_7542, n_7543, n_7544, n_7545;
  wire n_7546, n_7547, n_7548, n_7549, n_7550, n_7551, n_7552, n_7553;
  wire n_7554, n_7555, n_7556, n_7557, n_7558, n_7559, n_7560, n_7561;
  wire n_7562, n_7563, n_7564, n_7565, n_7566, n_7567, n_7568, n_7569;
  wire n_7570, n_7571, n_7572, n_7573, n_7574, n_7575, n_7576, n_7577;
  wire n_7578, n_7579, n_7580, n_7581, n_7582, n_7583, n_7584, n_7585;
  wire n_7586, n_7587, n_7588, n_7589, n_7590, n_7591, n_7592, n_7593;
  wire n_7596, n_7597, n_7598, n_7599, n_7600, n_7601, n_7602, n_7603;
  wire n_7604, n_7605, n_7606, n_7607, n_7608, n_7609, n_7610, n_7611;
  wire n_7612, n_7613, n_7614, n_7615, n_7616, n_7617, n_7618, n_7619;
  wire n_7620, n_7621, n_7622, n_7623, n_7624, n_7625, n_7626, n_7627;
  wire n_7628, n_7629, n_7630, n_7631, n_7632, n_7633, n_7635, n_7636;
  wire n_7669, n_7670, n_7671, n_7672, n_7673, n_7674, n_7675, n_7676;
  wire n_7677, n_7678, n_7680, n_7681, n_7682, n_7683, n_7684, n_7685;
  wire n_7686, n_7687, n_7688, n_7689, n_7690, n_7691, n_7692, n_7693;
  wire n_7694, n_7696, n_7697, n_7698, n_7699, n_7700, n_7701, n_7702;
  wire n_7703, n_7704, n_7705, n_7706, n_7707, n_7708, n_7709, n_7710;
  wire n_7711, n_7712, n_7713, n_7714, n_7715, n_7716, n_7717, n_7718;
  wire n_7719, n_7720, n_7721, n_7722, n_7723, n_7724, n_7725, n_7726;
  wire n_7727, n_7728, n_7729, n_7730, n_7731, n_7765, n_7766, n_7767;
  wire n_7768, n_7769, n_7770, n_7771, n_7772, n_7773, n_7774, n_7775;
  wire n_7776, n_7777, n_7778, n_7779, n_7780, n_7781, n_7782, n_7783;
  wire n_7784, n_7785, n_7786, n_7787, n_7788, n_7789, n_7790, n_7791;
  wire n_7792, n_7793, n_7794, n_7795, n_7796, n_7797, n_7798, n_7799;
  wire n_7800, n_7801, n_7802, n_7803, n_7804, n_7805, n_7806, n_7807;
  wire n_7808, n_7809, n_7810, n_7811, n_7812, n_7813, n_7814, n_7815;
  wire n_7816, n_7817, n_7818, n_7819, n_7820, n_7821, n_7822, n_7823;
  wire n_7824, n_7825, n_7827, n_7828, n_7829, n_7830, n_7831, n_7832;
  wire n_7833, n_7834, n_7835, n_7836, n_7837, n_7838, n_7839, n_7840;
  wire n_7841, n_7842, n_7843, n_7844, n_7845, n_7846, n_7847, n_7848;
  wire n_7849, n_7850, n_7851, n_7852, n_7853, n_7854, n_7855, n_7856;
  wire n_7857, n_7859, n_7860, n_7861, n_7862, n_7882, n_7883, n_7884;
  wire n_7885, n_7886, n_7887, n_7888, n_7889, n_7890, n_7891, n_7892;
  wire n_7893, n_7894, n_7895, n_7896, n_7897, n_7898, n_7899, n_7900;
  wire n_7901, n_7902, n_7903, n_7904, n_7905, n_7906, n_7907, n_7908;
  wire n_7909, n_7910, n_7911, n_7913, n_7914, n_7915, n_7916, n_7917;
  wire n_7918, n_7919, n_7921, n_7922, n_7923, n_7924, n_7925, n_7926;
  wire n_7927, n_7928, n_7929, n_7930, n_7931, n_7932, n_7933, n_7934;
  wire n_7935, n_7936, n_7937, n_7938, n_7939, n_7940, n_7941, n_7942;
  wire n_7943, n_7944, n_7945, n_7946, n_7947, n_7948, n_7949, n_7950;
  wire n_7951, n_7952, n_7953, n_7954, n_7955, n_7956, n_7957, n_7958;
  wire n_7959, n_7960, n_7961, n_7962, n_7963, n_7964, n_7965, n_7966;
  wire n_7967, n_7968, n_7969, n_7970, n_7971, n_7972, n_7973, n_7975;
  wire n_7976, n_7977, n_7978, n_7979, n_7980, n_7981, n_7982, n_7983;
  wire n_7984, n_7985, n_7986, n_7987, n_7988, n_7989, n_7990, n_7991;
  wire n_7992, n_7993, n_7994, n_7995, n_7996, n_7997, n_7998, n_7999;
  wire n_8000, n_8001, n_8002, n_8003, n_8004, n_8005, n_8006, n_8008;
  wire n_8009, n_8010, n_8011, n_8012, n_8013, n_8014, n_8015, n_8016;
  wire n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8024, n_8025;
  wire n_8026, n_8027, n_8028, n_8029, n_8030, n_8031, n_8032, n_8033;
  wire n_8034, n_8035, n_8036, n_8037, n_8038, n_8039, n_8040, n_8041;
  wire n_8042, n_8043, n_8044, n_8045, n_8046, n_8047, n_8048, n_8049;
  wire n_8050, n_8051, n_8052, n_8053, n_8054, n_8055, n_8056, n_8057;
  wire n_8058, n_8059, n_8060, n_8061, n_8062, n_8063, n_8064, n_8065;
  wire n_8066, n_8067, n_8068, n_8069, n_8070, n_8071, n_8072, n_8073;
  wire n_8074, n_8075, n_8076, n_8077, n_8078, n_8079, n_8080, n_8081;
  wire n_8082, n_8083, n_8084, n_8085, n_8086, n_8087, n_8088, n_8089;
  wire n_8090, n_8091, n_8092, n_8093, n_8094, n_8095, n_8096, n_8097;
  wire n_8098, n_8099, n_8100, n_8101, n_8102, n_8103, n_8104, n_8105;
  wire n_8106, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112, n_8113;
  wire n_8114, n_8115, n_8116, n_8117, n_8118, n_8119, n_8120, n_8121;
  wire n_8122, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128, n_8129;
  wire n_8130, n_8131, n_8132, n_8133, n_8134, n_8135, n_8136, n_8137;
  wire n_8138, n_8139, n_8140, n_8141, n_8142, n_8143, n_8144, n_8145;
  wire n_8146, n_8147, n_8148, n_8149, n_8150, n_8151, n_8152, n_8153;
  wire n_8154, n_8155, n_8156, n_8157, n_8158, n_8159, n_8160, n_8161;
  wire n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168, n_8169;
  wire n_8170, n_8171, n_8172, n_8173, n_8174, n_8175, n_8176, n_8177;
  wire n_8178, n_8179, n_8180, n_8181, n_8182, n_8183, n_8184, n_8185;
  wire n_8186, n_8187, n_8188, n_8189, n_8190, n_8191, n_8192, n_8193;
  wire n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200, n_8201;
  wire n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208, n_8209;
  wire n_8210, n_8211, n_8212, n_8213, n_8214, n_8215, n_8216, n_8217;
  wire n_8218, n_8219, n_8220, n_8221, n_8222, n_8223, n_8224, n_8225;
  wire n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232, n_8233;
  wire n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8240, n_8241;
  wire n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248, n_8249;
  wire n_8250, n_8251, n_8252, n_8253, n_8254, n_8255, n_8256, n_8257;
  wire n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264, n_8265;
  wire n_8266, n_8267, n_8268, n_8269, n_8270, n_8271, n_8272, n_8273;
  wire n_8274, n_8276, n_8280, n_8283, n_8284, n_8285, n_8286, n_8287;
  wire n_8288, n_8289, n_8292, n_8293, n_8294, n_8295, n_8296, n_8297;
  wire n_8300, n_8301, n_8302, n_8303, n_8304, n_8305, n_8306, n_8308;
  wire n_8309, n_8310, n_8311, n_8312, n_8313, n_8314, n_8315, n_8316;
  wire n_8317, n_8318, n_8320, n_8321, n_8322, n_8323, n_8326, n_8327;
  wire n_8329, n_8330, n_8331, n_8332, n_8333, n_8335, n_8337, n_8338;
  wire n_8339, n_8340, n_8341, n_8342, n_8343, n_8344, n_8345, n_8346;
  wire n_8347, n_8348, n_8349, n_8350, n_8351, n_8352, n_8353, n_8354;
  wire n_8355, n_8358, n_8359, n_8360, n_8361, n_8362, n_8363, n_8364;
  wire n_8365, n_8366, n_8370, n_8371, n_8372, n_8375, n_8376, n_8377;
  wire n_8378, n_8379, n_8382, n_8383, n_8386, n_8387, n_8388, n_8391;
  wire n_8392, n_8394, n_8396, n_8397, n_8398, n_8400, n_8401, n_8402;
  wire n_8403, n_8405, n_8411, n_8412, n_8413, n_8414, n_8415, n_8416;
  wire n_8417, n_8418, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424;
  wire n_8425, n_8426, n_8427, n_8428, n_8429, n_8430, n_8432, n_8433;
  wire n_8434, n_8435, n_8436, n_8438, n_8439, n_8440, n_8441, n_8442;
  wire n_8446, n_8450, n_8451, n_8453, n_8454, n_8456, n_8457, n_8458;
  wire n_8459, n_8460, n_8461, n_8462, n_8463, n_8464, n_8465, n_8467;
  wire n_8468, n_8469, n_8470, n_8471, n_8472, n_8473, n_8474, n_8475;
  wire n_8476, n_8477, n_8478, n_8479, n_8480, n_8481, n_8482, n_8484;
  wire n_8485, n_8486, n_8487, n_8488, n_8489, n_8490, n_8491, n_8492;
  wire n_8493, n_8494, n_8495, n_8496, n_8497, n_8499, n_8501, n_8502;
  wire n_8504, n_8505, n_8506, n_8508, n_8509, n_8510, n_8511, n_8512;
  wire n_8513, n_8514, n_8515, n_8516, n_8517, n_8518, n_8519, n_8520;
  wire n_8522, n_8523, n_8525, n_8526, n_8527, n_8528, n_8529, n_8530;
  wire n_8531, n_8532, n_8533, n_8534, n_8535, n_8536, n_8537, n_8538;
  wire n_8539, n_8540, n_8541, n_8542, n_8543, n_8544, n_8545, n_8546;
  wire n_8547, n_8548, n_8550, n_8551, n_8552, n_8553, n_8554, n_8555;
  wire n_8556, n_8557, n_8558, n_8559, n_8560, n_8561, n_8563, n_8564;
  wire n_8565, n_8566, n_8567, n_8568, n_8569, n_8570, n_8571, n_8576;
  wire n_8577, n_8578, n_8579, n_8587, n_8588, n_8589, n_8591, n_8592;
  wire n_8593, n_8594, n_8595, n_8596, n_8597, n_8598, n_8599, n_8600;
  wire n_8602, n_8603, n_8604, n_8605, n_8606, n_8607, n_8608, n_8609;
  wire n_8610, n_8611, n_8612, n_8613, n_8615, n_8616, n_8617, n_8618;
  wire n_8619, n_8620, n_8621, n_8622, n_8623, n_8624, n_8625, n_8652;
  wire n_8653, n_8654, n_8655, n_8656, n_8657, n_8658, n_8659, n_8660;
  wire n_8661, n_8662, n_8663, n_8664, n_8665, n_8666, n_8669, n_8670;
  wire n_8671, n_8673, n_8674, n_8675, n_8676, n_8677, n_8678, n_8680;
  wire n_8681, n_8682, n_8687, n_8688, n_8689, n_8690, n_8691, n_8692;
  wire n_8694, n_8695, n_8696, n_8697, n_8698, n_8699, n_8700, n_8701;
  wire n_8702, n_18079_BAR, n_18082_BAR, prev_load_request, rc_gclk,
       rc_gclk_199879, rc_gclk_199882, rc_gclk_199885;
  wire rc_gclk_199888, rc_gclk_199891, rc_gclk_199894, rc_gclk_199897,
       rc_gclk_199900, rc_gclk_199903, rc_gclk_199906, rc_gclk_199909;
  wire rc_gclk_199912, rc_gclk_199915, rc_gclk_199918, rc_gclk_199921,
       rc_gclk_199924, rc_gclk_199927, rc_gclk_199930, rc_gclk_199933;
  wire rc_gclk_199936, rc_gclk_199939, rc_gclk_199942, rc_gclk_199945,
       rc_gclk_199948, rc_gclk_199951, rc_gclk_199954, rc_gclk_199957;
  wire rc_gclk_199960, rc_gclk_199963, rc_gclk_199966, rc_gclk_199969,
       rc_gclk_199972, rc_gclk_199975, rc_gclk_199978, rc_gclk_199981;
  wire rc_gclk_199984, rc_gclk_199987, rc_gclk_199990, rc_gclk_199992,
       rc_gclk_199995, rc_gclk_199999, reset_internal_39074, reset_reg;
  wire \rs1_data[1]_39396 , \rs1_data[3]_39426 , \rs1_data[4]_39436 ,
       \rs1_data[6]_39456 , \rs1_data[7]_39466 , \rs1_data[9]_39486 ,
       \rs1_data[10]_39496 , \rs1_data[11]_39506 ;
  wire \rs1_data[12]_39516 , \rs1_data[13]_39536 , \rs1_data[14]_39546
       , \rs1_data[15]_39556 , \rs1_data[19]_39596 ,
       \rs1_data[21]_39616 , \rs1_data[22]_39626 , \rs1_data[23]_39326 ;
  wire \rs1_data[24]_39336 , \rs1_data[25]_39346 , \rs1_data[26]_39356
       , \rs1_data[29]_39416 , \rs1_data[30]_39526 , store_type,
       system_type, take_trap_39229;
  RC_CG_MOD_AUTO_rvsteel_core RC_CG_HIER_INST1(.ck_in (clock), .enable
       (n_8207), .test (1'b0), .ck_out (rc_gclk));
  RC_CG_MOD_AUTO_rvsteel_core_9 RC_CG_HIER_INST10(.ck_in (clock),
       .enable (n_8198), .test (1'b0), .ck_out (rc_gclk_199903));
  RC_CG_MOD_AUTO_rvsteel_core_10 RC_CG_HIER_INST11(.ck_in (clock),
       .enable (n_8197), .test (1'b0), .ck_out (rc_gclk_199906));
  RC_CG_MOD_AUTO_rvsteel_core_11 RC_CG_HIER_INST12(.ck_in (clock),
       .enable (n_8196), .test (1'b0), .ck_out (rc_gclk_199909));
  RC_CG_MOD_AUTO_rvsteel_core_12 RC_CG_HIER_INST13(.ck_in (clock),
       .enable (n_8195), .test (1'b0), .ck_out (rc_gclk_199912));
  RC_CG_MOD_AUTO_rvsteel_core_13 RC_CG_HIER_INST14(.ck_in (clock),
       .enable (n_8194), .test (1'b0), .ck_out (rc_gclk_199915));
  RC_CG_MOD_AUTO_rvsteel_core_14 RC_CG_HIER_INST15(.ck_in (clock),
       .enable (n_8193), .test (1'b0), .ck_out (rc_gclk_199918));
  RC_CG_MOD_AUTO_rvsteel_core_15 RC_CG_HIER_INST16(.ck_in (clock),
       .enable (n_8192), .test (1'b0), .ck_out (rc_gclk_199921));
  RC_CG_MOD_AUTO_rvsteel_core_16 RC_CG_HIER_INST17(.ck_in (clock),
       .enable (n_8191), .test (1'b0), .ck_out (rc_gclk_199924));
  RC_CG_MOD_AUTO_rvsteel_core_17 RC_CG_HIER_INST18(.ck_in (clock),
       .enable (n_8190), .test (1'b0), .ck_out (rc_gclk_199927));
  RC_CG_MOD_AUTO_rvsteel_core_18 RC_CG_HIER_INST19(.ck_in (clock),
       .enable (n_8189), .test (1'b0), .ck_out (rc_gclk_199930));
  RC_CG_MOD_AUTO_rvsteel_core_1 RC_CG_HIER_INST2(.ck_in (clock),
       .enable (n_8206), .test (1'b0), .ck_out (rc_gclk_199879));
  RC_CG_MOD_AUTO_rvsteel_core_19 RC_CG_HIER_INST20(.ck_in (clock),
       .enable (n_8188), .test (1'b0), .ck_out (rc_gclk_199933));
  RC_CG_MOD_AUTO_rvsteel_core_20 RC_CG_HIER_INST21(.ck_in (clock),
       .enable (n_8187), .test (1'b0), .ck_out (rc_gclk_199936));
  RC_CG_MOD_AUTO_rvsteel_core_21 RC_CG_HIER_INST22(.ck_in (clock),
       .enable (n_8186), .test (1'b0), .ck_out (rc_gclk_199939));
  RC_CG_MOD_AUTO_rvsteel_core_22 RC_CG_HIER_INST23(.ck_in (clock),
       .enable (n_8185), .test (1'b0), .ck_out (rc_gclk_199942));
  RC_CG_MOD_AUTO_rvsteel_core_23 RC_CG_HIER_INST24(.ck_in (clock),
       .enable (n_8184), .test (1'b0), .ck_out (rc_gclk_199945));
  RC_CG_MOD_AUTO_rvsteel_core_24 RC_CG_HIER_INST25(.ck_in (clock),
       .enable (n_8183), .test (1'b0), .ck_out (rc_gclk_199948));
  RC_CG_MOD_AUTO_rvsteel_core_25 RC_CG_HIER_INST26(.ck_in (clock),
       .enable (n_8182), .test (1'b0), .ck_out (rc_gclk_199951));
  RC_CG_MOD_AUTO_rvsteel_core_26 RC_CG_HIER_INST27(.ck_in (clock),
       .enable (n_8181), .test (1'b0), .ck_out (rc_gclk_199954));
  RC_CG_MOD_AUTO_rvsteel_core_27 RC_CG_HIER_INST28(.ck_in (clock),
       .enable (n_8180), .test (1'b0), .ck_out (rc_gclk_199957));
  RC_CG_MOD_AUTO_rvsteel_core_28 RC_CG_HIER_INST29(.ck_in (clock),
       .enable (n_8179), .test (1'b0), .ck_out (rc_gclk_199960));
  RC_CG_MOD_AUTO_rvsteel_core_2 RC_CG_HIER_INST3(.ck_in (clock),
       .enable (n_8205), .test (1'b0), .ck_out (rc_gclk_199882));
  RC_CG_MOD_AUTO_rvsteel_core_29 RC_CG_HIER_INST30(.ck_in (clock),
       .enable (n_8178), .test (1'b0), .ck_out (rc_gclk_199963));
  RC_CG_MOD_AUTO_rvsteel_core_30 RC_CG_HIER_INST31(.ck_in (clock),
       .enable (n_8177), .test (1'b0), .ck_out (rc_gclk_199966));
  RC_CG_MOD_AUTO_rvsteel_core_31 RC_CG_HIER_INST32(.ck_in (clock),
       .enable (n_8176), .test (1'b0), .ck_out (rc_gclk_199969));
  RC_CG_MOD_AUTO_rvsteel_core_32 RC_CG_HIER_INST33(.ck_in (clock),
       .enable (n_8175), .test (1'b0), .ck_out (rc_gclk_199972));
  RC_CG_MOD_AUTO_rvsteel_core_33 RC_CG_HIER_INST34(.ck_in (clock),
       .enable (n_8174), .test (1'b0), .ck_out (rc_gclk_199975));
  RC_CG_MOD_AUTO_rvsteel_core_34 RC_CG_HIER_INST35(.ck_in (clock),
       .enable (n_8173), .test (1'b0), .ck_out (rc_gclk_199978));
  RC_CG_MOD_AUTO_rvsteel_core_35 RC_CG_HIER_INST36(.ck_in (clock),
       .enable (n_8172), .test (1'b0), .ck_out (rc_gclk_199981));
  RC_CG_MOD_AUTO_rvsteel_core_36 RC_CG_HIER_INST37(.ck_in (clock),
       .enable (n_8171), .test (1'b0), .ck_out (rc_gclk_199984));
  RC_CG_MOD_AUTO_rvsteel_core_37 RC_CG_HIER_INST38(.ck_in (clock),
       .enable (n_8170), .test (1'b0), .ck_out (rc_gclk_199987));
  RC_CG_MOD_AUTO_rvsteel_core_38 RC_CG_HIER_INST39(.ck_in (clock),
       .enable (n_8169), .test (1'b0), .ck_out (rc_gclk_199990));
  RC_CG_MOD_AUTO_rvsteel_core_3 RC_CG_HIER_INST4(.ck_in (clock),
       .enable (n_8204), .test (1'b0), .ck_out (rc_gclk_199885));
  RC_CG_MOD_AUTO_rvsteel_core_39 RC_CG_HIER_INST40(.ck_in (clock),
       .enable (n_7305), .test (1'b0), .ck_out (rc_gclk_199992));
  RC_CG_MOD_AUTO_rvsteel_core_40 RC_CG_HIER_INST41(.ck_in (clock),
       .enable (n_8168), .test (1'b0), .ck_out (rc_gclk_199995));
  RC_CG_MOD_AUTO_rvsteel_core_41 RC_CG_HIER_INST42(.ck_in (clock),
       .enable (n_8167), .test (1'b0), .ck_out (rc_gclk_199999));
  RC_CG_MOD_AUTO_rvsteel_core_4 RC_CG_HIER_INST5(.ck_in (clock),
       .enable (n_8203), .test (1'b0), .ck_out (rc_gclk_199888));
  RC_CG_MOD_AUTO_rvsteel_core_5 RC_CG_HIER_INST6(.ck_in (clock),
       .enable (n_8202), .test (1'b0), .ck_out (rc_gclk_199891));
  RC_CG_MOD_AUTO_rvsteel_core_6 RC_CG_HIER_INST7(.ck_in (clock),
       .enable (n_8201), .test (1'b0), .ck_out (rc_gclk_199894));
  RC_CG_MOD_AUTO_rvsteel_core_7 RC_CG_HIER_INST8(.ck_in (clock),
       .enable (n_8200), .test (1'b0), .ck_out (rc_gclk_199897));
  RC_CG_MOD_AUTO_rvsteel_core_8 RC_CG_HIER_INST9(.ck_in (clock),
       .enable (n_8199), .test (1'b0), .ck_out (rc_gclk_199900));
  csa_tree_add_1660_20_group_293 csa_tree_add_1660_20_groupi(.in_0
       ({n_6134, \rs1_data[30]_39526 , \rs1_data[29]_39416 , n_6136,
       n_6135, n_6161, \rs1_data[25]_39346 , n_6145, n_6143, n_6159,
       \rs1_data[21]_39616 , n_6149, \rs1_data[19]_39596 , n_6141,
       n_8366, n_6132, n_6155, n_6153, \rs1_data[13]_39536 ,
       \rs1_data[12]_39516 , \rs1_data[11]_39506 , n_6139, n_6137,
       n_6127, n_6183, n_6165, n_6170, n_6178, n_6181, n_6123, n_6167,
       n_6121}), .in_1 ({UNCONNECTED_HIER_Z0, UNCONNECTED_HIER_Z,
       n_8264, n_8265, n_8266, n_8267, n_8268, n_8269, n_8270, n_8271,
       n_8272, n_8273, n_8274, n_8491, n_8276, n_8314, n_8312, n_8315,
       n_8280, n_8490, n_8311, n_8283, n_8284, n_8285, n_8286, n_8287,
       n_8288, n_8289, n_8313, n_8316, n_8292, n_8293, n_8294,
       n_8295}), .in_2 ({UNCONNECTED_HIER_Z33, UNCONNECTED_HIER_Z32,
       UNCONNECTED_HIER_Z31, UNCONNECTED_HIER_Z30,
       UNCONNECTED_HIER_Z29, UNCONNECTED_HIER_Z28,
       UNCONNECTED_HIER_Z27, UNCONNECTED_HIER_Z26,
       UNCONNECTED_HIER_Z25, UNCONNECTED_HIER_Z24,
       UNCONNECTED_HIER_Z23, UNCONNECTED_HIER_Z22,
       UNCONNECTED_HIER_Z21, UNCONNECTED_HIER_Z20,
       UNCONNECTED_HIER_Z19, UNCONNECTED_HIER_Z18,
       UNCONNECTED_HIER_Z17, UNCONNECTED_HIER_Z16,
       UNCONNECTED_HIER_Z15, UNCONNECTED_HIER_Z14,
       UNCONNECTED_HIER_Z13, UNCONNECTED_HIER_Z12,
       UNCONNECTED_HIER_Z11, UNCONNECTED_HIER_Z10, UNCONNECTED_HIER_Z9,
       UNCONNECTED_HIER_Z8, UNCONNECTED_HIER_Z7, UNCONNECTED_HIER_Z6,
       UNCONNECTED_HIER_Z5, UNCONNECTED_HIER_Z4, UNCONNECTED_HIER_Z3,
       UNCONNECTED_HIER_Z2, UNCONNECTED_HIER_Z1,
       alu_operation_code_39112}), .out_0 ({n_7696, n_7697, n_7698,
       n_7699, n_7700, n_7701, n_7702, n_7703, n_7704, n_7705, n_7706,
       n_7709, n_7711, n_7712, n_7713, n_7715, n_7716, n_7717, n_7718,
       n_7719, n_7720, n_7721, n_7722, n_7723, n_7724, n_7725, n_7726,
       n_7727, n_7728, n_7729, n_7730, n_7731}));
  BUX1 g27809(.A (n_7627), .Q (rw_address[31]));
  BUX1 g27788(.A (n_7601), .Q (rw_address[17]));
  BUX1 g27803(.A (n_7597), .Q (rw_address[21]));
  BUX1 g27792(.A (n_7622), .Q (rw_address[25]));
  BUX1 g27800(.A (n_7617), .Q (rw_address[29]));
  BUX1 g27812(.A (n_7624), .Q (rw_address[23]));
  BUX1 g27805(.A (n_7620), .Q (rw_address[27]));
  BUX1 g27810(.A (n_7606), .Q (rw_address[30]));
  BUX1 g27799(.A (n_7621), .Q (rw_address[26]));
  BUX1 g27795(.A (n_7599), .Q (rw_address[19]));
  BUX1 g27815(.A (n_7619), .Q (rw_address[28]));
  BUX1 g27806(.A (n_7596), .Q (rw_address[22]));
  BUX1 g27791(.A (n_7600), .Q (rw_address[18]));
  BUX1 g27798(.A (n_7598), .Q (rw_address[20]));
  BUX1 g27816(.A (n_7602), .Q (rw_address[16]));
  BUX1 g27796(.A (n_7612), .Q (rw_address[7]));
  BUX1 g27811(.A (n_7604), .Q (rw_address[14]));
  BUX1 g27808(.A (n_7605), .Q (rw_address[13]));
  BUX1 g27807(.A (n_7607), .Q (rw_address[12]));
  BUX1 g27801(.A (n_7610), .Q (rw_address[9]));
  BUX1 g27802(.A (n_7609), .Q (rw_address[10]));
  BUX1 g27797(.A (n_7611), .Q (rw_address[8]));
  BUX1 g27794(.A (n_7613), .Q (rw_address[6]));
  BUX1 g27793(.A (n_7614), .Q (rw_address[5]));
  BUX1 g27790(.A (n_7615), .Q (rw_address[4]));
  BUX1 g27789(.A (n_7616), .Q (rw_address[3]));
  BUX1 g27814(.A (n_7623), .Q (rw_address[24]));
  BUX1 g27804(.A (n_7608), .Q (rw_address[11]));
  BUX1 g27787(.A (n_7618), .Q (rw_address[2]));
  BUX1 g27785(.A (n_7625), .Q (rw_address[0]));
  BUX1 g27813(.A (n_7603), .Q (rw_address[15]));
  BUX1 g27784(.A (n_7626), .Q (rw_address[1]));
  BUX1 g27786(.A (n_7630), .Q (write_strobe[0]));
  BUX1 g27783(.A (n_7628), .Q (write_strobe[3]));
  BUX1 g27782(.A (n_7631), .Q (write_strobe[2]));
  BUX1 g27781(.A (n_7629), .Q (write_strobe[1]));
  INX1 g27817(.A (n_8160), .Q (n_6195));
  BUX2 g27825(.A (n_7400), .Q (n_6237));
  BUX1 g27822(.A (n_7399), .Q (n_6238));
  BUX3 g27839(.A (n_8208), .Q (n_6234));
  BUX2 g27828(.A (n_7633), .Q (n_6233));
  BUX2 g27833(.A (n_7401), .Q (n_6232));
  BUX2 g27830(.A (n_7636), .Q (n_6236));
  BUX1 g27884(.A (n_6126), .Q (n_6165));
  BUX1 g27911(.A (\rs1_data[3]_39426 ), .Q (n_6181));
  BUX1 g27893(.A (\rs1_data[4]_39436 ), .Q (n_6178));
  BUX1 g27908(.A (n_2306), .Q (n_6170));
  BUX1 g27915(.A (\rs1_data[1]_39396 ), .Q (n_6167));
  BUX1 g27880(.A (\rs1_data[7]_39466 ), .Q (n_6183));
  BUX2 g27843(.A (alu_sra_result[31]), .Q (n_6134));
  BUX1 g27854(.A (\rs1_data[26]_39356 ), .Q (n_6161));
  BUX1 g27863(.A (\rs1_data[15]_39556 ), .Q (n_6155));
  BUX1 g27860(.A (\rs1_data[22]_39626 ), .Q (n_6159));
  BUX1 g27866(.A (\rs1_data[14]_39546 ), .Q (n_6153));
  BUX1 g27868(.A (\rs1_data[24]_39336 ), .Q (n_6145));
  BUX1 g27857(.A (\rs1_data[23]_39326 ), .Q (n_6143));
  BUX1 g27877(.A (\rs1_data[10]_39496 ), .Q (n_6139));
  BUX1 g27905(.A (\rs1_data[9]_39486 ), .Q (n_6137));
  BUX1 g27885(.A (\rs1_data[6]_39456 ), .Q (n_6126));
  INX1 g27929(.A (prev_rw_address[27]), .Q (n_6114));
  INX1 g27920(.A (prev_rw_address[28]), .Q (n_6113));
  INX1 g27922(.A (prev_rw_address[29]), .Q (n_6112));
  INX1 g27919(.A (prev_rw_address[2]), .Q (n_6111));
  INX1 g27938(.A (prev_rw_address[30]), .Q (n_6110));
  INX1 g27921(.A (prev_rw_address[31]), .Q (n_6109));
  INX1 g27923(.A (prev_rw_address[3]), .Q (n_6108));
  INX1 g27933(.A (prev_rw_address[4]), .Q (n_6107));
  INX1 g27934(.A (prev_rw_address[5]), .Q (n_6106));
  INX1 g27928(.A (prev_rw_address[6]), .Q (n_6105));
  INX1 g27925(.A (prev_rw_address[7]), .Q (n_6104));
  INX1 g27927(.A (prev_rw_address[8]), .Q (n_6103));
  INX1 g27937(.A (prev_rw_address[9]), .Q (n_6102));
  INX1 g27943(.A (prev_rw_address[10]), .Q (n_6101));
  INX1 g27940(.A (prev_rw_address[11]), .Q (n_6100));
  INX1 g27931(.A (prev_rw_address[12]), .Q (n_6099));
  INX1 g27947(.A (prev_rw_address[13]), .Q (n_6098));
  INX1 g27944(.A (prev_rw_address[14]), .Q (n_6097));
  INX1 g27945(.A (prev_rw_address[15]), .Q (n_6096));
  INX1 g27924(.A (prev_rw_address[16]), .Q (n_6095));
  INX1 g27946(.A (prev_rw_address[17]), .Q (n_6094));
  INX1 g27926(.A (prev_rw_address[18]), .Q (n_6093));
  INX1 g27941(.A (prev_rw_address[19]), .Q (n_6092));
  INX1 g27942(.A (prev_rw_address[20]), .Q (n_6091));
  INX1 g27930(.A (prev_rw_address[21]), .Q (n_6090));
  INX1 g27948(.A (prev_rw_address[22]), .Q (n_6089));
  INX1 g27932(.A (prev_rw_address[23]), .Q (n_6088));
  INX1 g27939(.A (prev_rw_address[24]), .Q (n_6087));
  INX1 g27935(.A (prev_rw_address[25]), .Q (n_6086));
  INX1 g27936(.A (prev_rw_address[26]), .Q (n_6085));
  INX1 g27949(.A (csr_mscratch[2]), .Q (n_6084));
  INX1 g27952(.A (prev_instruction[18]), .Q (n_6083));
  BUX1 g27953(.A (current_state[2]), .Q (n_6082));
  NA3X4 g50684(.A (n_8615), .B (n_6052), .C (n_6049), .Q (n_6121));
  NA3I1X4 g50685(.B (n_5961), .C (n_6072), .AN (n_6047), .Q (n_6136));
  NA3X4 g50686(.A (n_5955), .B (n_6079), .C (n_6043), .Q
       (\rs1_data[15]_39556 ));
  NA3X4 g50687(.A (n_8400), .B (n_8624), .C (n_6040), .Q
       (\rs1_data[13]_39536 ));
  NA3X4 g50688(.A (n_5958), .B (n_6066), .C (n_6045), .Q
       (\rs1_data[30]_39526 ));
  NA3X4 g50689(.A (n_8401), .B (n_8602), .C (n_8604), .Q
       (\rs1_data[21]_39616 ));
  NA3X4 g50690(.A (n_8610), .B (n_6075), .C (n_6034), .Q
       (\rs1_data[23]_39326 ));
  NA3X4 g50691(.A (n_8398), .B (n_6074), .C (n_6035), .Q
       (\rs1_data[24]_39336 ));
  NA3X2 g50692(.A (n_5956), .B (n_6077), .C (n_6046), .Q
       (\rs1_data[26]_39356 ));
  NA3I1X4 g50693(.B (n_8397), .C (n_6073), .AN (n_6044), .Q
       (alu_sra_result[31]));
  NA3X4 g50694(.A (n_5957), .B (n_6078), .C (n_6041), .Q
       (\rs1_data[10]_39496 ));
  NA3X4 g50695(.A (n_5947), .B (n_6076), .C (n_6036), .Q
       (\rs1_data[29]_39416 ));
  NA3I1X2 g50696(.B (n_5962), .C (n_4525), .AN (n_6027), .Q
       (\rs1_data[22]_39626 ));
  NA3I1X4 g50697(.B (n_5959), .C (n_6071), .AN (n_6042), .Q
       (\rs1_data[14]_39546 ));
  NA3X4 g50698(.A (n_5951), .B (n_6064), .C (n_6038), .Q
       (\rs1_data[12]_39516 ));
  NA3I1X4 g50699(.B (n_8405), .C (n_6065), .AN (n_6025), .Q
       (\rs1_data[25]_39346 ));
  NA3X4 g50700(.A (n_5935), .B (n_6054), .C (n_5975), .Q (n_2306));
  NA3X4 g50701(.A (n_5945), .B (n_6068), .C (n_6033), .Q (n_6135));
  NA3X4 g50702(.A (n_5941), .B (n_6062), .C (n_6023), .Q (n_6132));
  NA3I1X4 g50703(.B (n_5950), .C (n_6080), .AN (n_6037), .Q
       (\rs1_data[11]_39506 ));
  NA3X4 g50704(.A (n_5942), .B (n_6067), .C (n_6039), .Q (n_6149));
  NA3I1X4 g50705(.B (n_8402), .C (n_6061), .AN (n_6024), .Q (n_6141));
  NA3I1X4 g50706(.B (n_8611), .C (n_8603), .AN (n_6012), .Q
       (\rs1_data[9]_39486 ));
  NA3I1X4 g50708(.B (n_8612), .C (n_6056), .AN (n_5990), .Q
       (\rs1_data[6]_39456 ));
  NA3X4 g50709(.A (n_5938), .B (n_6058), .C (n_5998), .Q (n_6127));
  NA3X4 g50710(.A (n_8613), .B (n_6057), .C (n_8694), .Q
       (\rs1_data[7]_39466 ));
  NA3I1X4 g50711(.B (n_5936), .C (n_6055), .AN (n_5989), .Q
       (\rs1_data[3]_39426 ));
  NA3X4 g50712(.A (n_6053), .B (n_5933), .C (n_5976), .Q (n_6123));
  NA3I1X4 g50713(.B (n_8625), .C (n_8370), .AN (n_8391), .Q
       (\rs1_data[4]_39436 ));
  NA3X4 g50714(.A (n_5932), .B (n_6050), .C (n_5972), .Q
       (\rs1_data[1]_39396 ));
  NA3X4 g50715(.A (n_8403), .B (n_6070), .C (n_6028), .Q
       (\rs1_data[19]_39596 ));
  NO2X2 g50716(.A (n_6011), .B (n_8607), .Q (n_6080));
  NO2X2 g50717(.A (n_8372), .B (n_6013), .Q (n_6079));
  NO2X2 g50718(.A (n_8605), .B (n_8377), .Q (n_6078));
  NO2X2 g50719(.A (n_6017), .B (n_6015), .Q (n_6077));
  NO2X2 g50720(.A (n_6026), .B (n_6009), .Q (n_6076));
  NO2X2 g50721(.A (n_8376), .B (n_5984), .Q (n_6075));
  NO2X2 g50722(.A (n_6048), .B (n_6000), .Q (n_6074));
  AND6X2 g50726(.A (n_8415), .B (n_8424), .C (n_5716), .D (n_5724), .E
       (n_5695), .F (n_5798), .Q (n_6071));
  NO2X2 g50727(.A (n_8382), .B (n_6007), .Q (n_6070));
  NO2X2 g50729(.A (n_6008), .B (n_6006), .Q (n_6068));
  NO2X2 g50730(.A (n_6003), .B (n_5996), .Q (n_6067));
  NO2X2 g50731(.A (n_8371), .B (n_8378), .Q (n_6066));
  NO2X2 g50732(.A (n_8379), .B (n_8383), .Q (n_6065));
  NO2X2 g50733(.A (n_6022), .B (n_5994), .Q (n_6064));
  NO2X4 g50735(.A (n_8375), .B (n_5991), .Q (n_6062));
  NO3X2 g50736(.A (n_5992), .B (n_5892), .C (n_5893), .Q (n_6061));
  NO2X2 g50737(.A (n_8386), .B (n_5986), .Q (n_6060));
  NO2X2 g50739(.A (n_8606), .B (n_5980), .Q (n_6058));
  NO2X2 g50740(.A (n_8387), .B (n_5979), .Q (n_6057));
  NO2X2 g50741(.A (n_8388), .B (n_5978), .Q (n_6056));
  NO2X4 g50742(.A (n_8608), .B (n_8695), .Q (n_6055));
  NO3X4 g50743(.A (n_8392), .B (n_5806), .C (n_5816), .Q (n_6054));
  NO2X4 g50744(.A (n_8609), .B (n_5973), .Q (n_6053));
  NO2X4 g50745(.A (n_8394), .B (n_5965), .Q (n_6052));
  NO2X2 g50747(.A (n_8396), .B (n_5964), .Q (n_6050));
  NO2X2 g50748(.A (n_5340), .B (n_5963), .Q (n_6049));
  NA3X1 g50749(.A (n_8421), .B (n_5694), .C (n_5624), .Q (n_6048));
  NA3X1 g50750(.A (n_5399), .B (n_5887), .C (n_5734), .Q (n_6047));
  AND4X1 g50751(.A (n_5398), .B (n_5681), .C (n_5688), .D (n_5574), .Q
       (n_6046));
  AND3X1 g50752(.A (n_5395), .B (n_8435), .C (n_5686), .Q (n_6045));
  NA3X1 g50753(.A (n_5400), .B (n_5927), .C (n_5594), .Q (n_6044));
  AND3X1 g50754(.A (n_5397), .B (n_8417), .C (n_5573), .Q (n_6043));
  NA3X1 g50755(.A (n_5396), .B (n_8412), .C (n_5593), .Q (n_6042));
  AND3X1 g50756(.A (n_5886), .B (n_5380), .C (n_5683), .Q (n_6041));
  NO2X1 g50757(.A (n_5930), .B (n_5858), .Q (n_6040));
  AND3X1 g50758(.A (n_5375), .B (n_5857), .C (n_5600), .Q (n_6039));
  AND3X1 g50759(.A (n_5377), .B (n_5875), .C (n_5531), .Q (n_6038));
  NA3X1 g50760(.A (n_5376), .B (n_8436), .C (n_5530), .Q (n_6037));
  AND3X1 g50761(.A (n_5379), .B (n_8441), .C (n_5672), .Q (n_6036));
  AND3X1 g50762(.A (n_5382), .B (n_8438), .C (n_5630), .Q (n_6035));
  AND3X1 g50763(.A (n_5381), .B (n_8439), .C (n_5629), .Q (n_6034));
  AND3X2 g50764(.A (n_5378), .B (n_5863), .C (n_5626), .Q (n_6033));
  AND3X1 g50769(.A (n_5374), .B (n_8670), .C (n_5669), .Q (n_6028));
  NA3X1 g50770(.A (n_5401), .B (n_8669), .C (n_5735), .Q (n_6027));
  NA3X1 g50771(.A (n_8422), .B (n_5692), .C (n_5620), .Q (n_6026));
  NA3X1 g50772(.A (n_5373), .B (n_8442), .C (n_5604), .Q (n_6025));
  NA3X1 g50773(.A (n_5856), .B (n_5368), .C (n_5599), .Q (n_6024));
  AND3X1 g50774(.A (n_5855), .B (n_5367), .C (n_5598), .Q (n_6023));
  NA2X1 g50775(.A (n_8426), .B (n_5885), .Q (n_6022));
  NA3X1 g50780(.A (n_8411), .B (n_5730), .C (n_5666), .Q (n_6017));
  NA2X1 g50782(.A (n_8419), .B (n_5862), .Q (n_6015));
  NA2X1 g50784(.A (n_5911), .B (n_8440), .Q (n_6013));
  NA3X1 g50785(.A (n_5350), .B (n_8446), .C (n_5514), .Q (n_6012));
  NA2X1 g50786(.A (n_8428), .B (n_8427), .Q (n_6011));
  NA3X1 g50788(.A (n_5881), .B (n_5566), .C (n_5572), .Q (n_6009));
  NA3X1 g50789(.A (n_5879), .B (n_5570), .C (n_5564), .Q (n_6008));
  NA3X1 g50790(.A (n_8423), .B (n_5619), .C (n_5618), .Q (n_6007));
  NA3X2 g50791(.A (n_5907), .B (n_5617), .C (n_5616), .Q (n_6006));
  NA2X1 g50794(.A (n_5870), .B (n_5851), .Q (n_6003));
  NA3X1 g50797(.A (n_5877), .B (n_5547), .C (n_5560), .Q (n_6000));
  NO2X2 g50799(.A (n_5906), .B (n_5828), .Q (n_5998));
  NA3X1 g50801(.A (n_8430), .B (n_5585), .C (n_5584), .Q (n_5996));
  NO2X1 g50802(.A (n_5919), .B (n_5837), .Q (n_5995));
  NA2X1 g50803(.A (n_5873), .B (n_5845), .Q (n_5994));
  NA2X1 g50805(.A (n_5869), .B (n_5843), .Q (n_5992));
  NA2X1 g50806(.A (n_5868), .B (n_5842), .Q (n_5991));
  NA3X1 g50807(.A (n_5346), .B (n_5826), .C (n_5502), .Q (n_5990));
  NA3X1 g50808(.A (n_5341), .B (n_5825), .C (n_5465), .Q (n_5989));
  NA2X1 g50811(.A (n_5840), .B (n_5831), .Q (n_5986));
  NA3X1 g50813(.A (n_5880), .B (n_5552), .C (n_5558), .Q (n_5984));
  NA3X2 g50817(.A (n_5822), .B (n_4792), .C (n_5520), .Q (n_5980));
  NA3X1 g50818(.A (n_5821), .B (n_4791), .C (n_5518), .Q (n_5979));
  NA3X1 g50819(.A (n_5820), .B (n_4790), .C (n_5516), .Q (n_5978));
  NO2X2 g50821(.A (n_5819), .B (n_5803), .Q (n_5976));
  NO2X2 g50822(.A (n_5824), .B (n_5815), .Q (n_5975));
  NA3X2 g50824(.A (n_8702), .B (n_5461), .C (n_5463), .Q (n_5973));
  NO3X2 g50825(.A (n_8698), .B (n_5453), .C (n_8464), .Q (n_5972));
  NA2X4 g50832(.A (n_5804), .B (n_5801), .Q (n_5965));
  NA3X2 g50833(.A (n_5799), .B (n_5460), .C (n_5422), .Q (n_5964));
  NA3X2 g50834(.A (n_5444), .B (n_5608), .C (n_5421), .Q (n_5963));
  NO2X1 g50835(.A (n_5795), .B (n_5796), .Q (n_5962));
  AND4X1 g50836(.A (n_5412), .B (n_5413), .C (n_5416), .D (n_5326), .Q
       (n_5961));
  NO2X1 g50838(.A (n_5797), .B (n_5793), .Q (n_5959));
  NO2X1 g50839(.A (n_5791), .B (n_5792), .Q (n_5958));
  NO2X1 g50840(.A (n_5787), .B (n_5790), .Q (n_5957));
  NO2X1 g50841(.A (n_5786), .B (n_5789), .Q (n_5956));
  NO2X1 g50842(.A (n_5785), .B (n_5788), .Q (n_5955));
  NO2X2 g50846(.A (n_5766), .B (n_5767), .Q (n_5951));
  NO2X1 g50847(.A (n_5764), .B (n_5765), .Q (n_5950));
  NO2X1 g50850(.A (n_5776), .B (n_5777), .Q (n_5947));
  NO2X1 g50852(.A (n_5772), .B (n_5773), .Q (n_5945));
  NO2X1 g50855(.A (n_5782), .B (n_5771), .Q (n_5942));
  NO2X1 g50856(.A (n_5781), .B (n_5770), .Q (n_5941));
  NO2X2 g50859(.A (n_5756), .B (n_8699), .Q (n_5938));
  NO2X2 g50861(.A (n_8454), .B (n_5754), .Q (n_5936));
  NO2X1 g50862(.A (n_5747), .B (n_5748), .Q (n_5935));
  NO2X4 g50864(.A (n_5741), .B (n_5745), .Q (n_5933));
  NO3X2 g50865(.A (n_5744), .B (n_8675), .C (n_8478), .Q (n_5932));
  NA3X1 g50867(.A (n_5603), .B (n_4828), .C (n_4827), .Q (n_5930));
  NA2X4 g50869(.A (n_5736), .B (n_4715), .Q (n_7682));
  NA2X4 g50870(.A (n_5739), .B (n_4716), .Q (n_7680));
  NA2X4 g50871(.A (n_5737), .B (n_4714), .Q (n_7681));
  NA2X2 g50872(.A (n_5738), .B (n_4713), .Q (n_2437));
  AND2X1 g50874(.A (n_5708), .B (n_5733), .Q (n_5927));
  AN21X1 g50877(.A (n_4741), .B (n_7187), .C (n_5702), .Q (n_5924));
  NA2X1 g50882(.A (n_5349), .B (n_5500), .Q (n_5919));
  NO2X1 g50891(.A (n_4996), .B (n_5680), .Q (n_5911));
  NO2X1 g50895(.A (n_5690), .B (n_5670), .Q (n_5907));
  NA2X1 g50896(.A (n_8477), .B (n_5512), .Q (n_5906));
  AND2X1 g50899(.A (n_5613), .B (n_5633), .Q (n_5904));
  AND2X1 g50900(.A (n_5614), .B (n_5632), .Q (n_5903));
  NA2X1 g50910(.A (n_5645), .B (n_5583), .Q (n_5893));
  NA2X1 g50911(.A (n_5653), .B (n_5582), .Q (n_5892));
  AND2X1 g50916(.A (n_5709), .B (n_5595), .Q (n_5887));
  NO2X1 g50917(.A (n_5689), .B (n_5575), .Q (n_5886));
  NO2X2 g50918(.A (n_5591), .B (n_5657), .Q (n_5885));
  NO2X1 g50919(.A (n_8673), .B (n_5655), .Q (n_5884));
  NO2X1 g50922(.A (n_4852), .B (n_5662), .Q (n_5881));
  NO2X1 g50923(.A (n_4853), .B (n_5663), .Q (n_5880));
  NO2X1 g50924(.A (n_4851), .B (n_5661), .Q (n_5879));
  AN21X1 g50925(.A (n_4741), .B (n_7094), .C (n_5660), .Q (n_5878));
  NO2X1 g50926(.A (n_4850), .B (n_5659), .Q (n_5877));
  NO2X1 g50928(.A (n_5610), .B (n_5602), .Q (n_5875));
  NO2X1 g50930(.A (n_4849), .B (n_5642), .Q (n_5873));
  NO2X1 g50932(.A (n_4847), .B (n_5640), .Q (n_5871));
  NO2X1 g50933(.A (n_4846), .B (n_5639), .Q (n_5870));
  NO2X1 g50934(.A (n_4845), .B (n_5638), .Q (n_5869));
  NO2X1 g50935(.A (n_4844), .B (n_5637), .Q (n_5868));
  NO2X1 g50940(.A (n_5668), .B (n_5542), .Q (n_5863));
  NO2X1 g50942(.A (n_5569), .B (n_5563), .Q (n_5862));
  NA2X1 g50947(.A (n_5611), .B (n_5532), .Q (n_5858));
  NO2X1 g50948(.A (n_5607), .B (n_5527), .Q (n_5857));
  NO2X1 g50949(.A (n_5606), .B (n_5526), .Q (n_5856));
  NO2X1 g50950(.A (n_5605), .B (n_5524), .Q (n_5855));
  NO2X1 g50954(.A (n_5557), .B (n_5551), .Q (n_5851));
  NO2X2 g50957(.A (n_5554), .B (n_5548), .Q (n_5848));
  NO2X1 g50959(.A (n_5540), .B (n_5536), .Q (n_5847));
  AND3X1 g50961(.A (n_5493), .B (n_5198), .C (n_5197), .Q (n_5845));
  NO2X1 g50963(.A (n_5522), .B (n_5491), .Q (n_5843));
  NO2X1 g50964(.A (n_5521), .B (n_5490), .Q (n_5842));
  NO2X1 g50965(.A (n_4824), .B (n_5534), .Q (n_5841));
  NO2X1 g50966(.A (n_4823), .B (n_5533), .Q (n_5840));
  NA2X1 g50971(.A (n_5505), .B (n_5507), .Q (n_5837));
  NO2X1 g50977(.A (n_5485), .B (n_5483), .Q (n_5831));
  NA2X1 g50982(.A (n_5715), .B (n_5228), .Q (n_7690));
  AO21X2 g50983(.A (n_8479), .B (n_8487), .C (n_5229), .Q (n_7689));
  AO21X1 g50984(.A (n_8479), .B (n_4640), .C (n_5229), .Q (n_7683));
  AO21X2 g50985(.A (n_8479), .B (n_4643), .C (n_5229), .Q (n_7686));
  AO21X1 g50986(.A (n_8479), .B (instruction[18]), .C (n_5229), .Q
       (n_7684));
  AO21X2 g50987(.A (n_8479), .B (instruction[17]), .C (n_5229), .Q
       (n_7685));
  NA2X1 g50988(.A (n_5504), .B (n_5489), .Q (n_5828));
  NO2X1 g50990(.A (n_5487), .B (n_5508), .Q (n_5826));
  NO2X2 g50991(.A (n_5475), .B (n_8459), .Q (n_5825));
  ON21X4 g50992(.A (n_5228), .B (branch_type), .C (n_4710), .Q
       (n_7691));
  NA3X1 g50993(.A (n_4765), .B (n_4766), .C (n_8618), .Q (n_5824));
  AND3X2 g50994(.A (n_4763), .B (n_4764), .C (n_5427), .Q (n_5823));
  AND2X1 g50995(.A (n_5474), .B (n_5478), .Q (n_5822));
  NO2X1 g50996(.A (n_8460), .B (n_5477), .Q (n_5821));
  NO2X1 g50997(.A (n_5472), .B (n_5476), .Q (n_5820));
  NA3X2 g50998(.A (n_4761), .B (n_4762), .C (n_5431), .Q (n_5819));
  NA2X1 g51001(.A (n_5462), .B (n_5464), .Q (n_5816));
  NA2X1 g51002(.A (n_8463), .B (n_8465), .Q (n_5815));
  AND2X1 g51010(.A (n_5440), .B (n_5449), .Q (n_5808));
  NA2X1 g51013(.A (n_4781), .B (n_5459), .Q (n_5806));
  NO3X2 g51016(.A (n_4778), .B (n_4510), .C (n_4511), .Q (n_5805));
  AND2X4 g51017(.A (n_4777), .B (n_5452), .Q (n_5804));
  NA2X1 g51018(.A (n_5466), .B (n_5426), .Q (n_5803));
  NO2X2 g51020(.A (n_8674), .B (n_5424), .Q (n_5801));
  NO3X1 g51022(.A (n_5121), .B (n_5045), .C (n_4717), .Q (n_5799));
  AN22X1 g51023(.A (n_4452), .B (n_6964), .C (n_4882), .D (n_6965), .Q
       (n_5798));
  OR4X1 g51024(.A (n_5018), .B (n_5020), .C (n_5019), .D (n_5021), .Q
       (n_5797));
  OR4X1 g51025(.A (n_5026), .B (n_5027), .C (n_4973), .D (n_5037), .Q
       (n_5796));
  OR4X1 g51026(.A (n_5024), .B (n_5035), .C (n_5025), .D (n_5036), .Q
       (n_5795));
  OR4X1 g51028(.A (n_5028), .B (n_5029), .C (n_5030), .D (n_5031), .Q
       (n_5793));
  OR4X1 g51029(.A (n_5005), .B (n_5006), .C (n_5017), .D (n_5016), .Q
       (n_5792));
  OR4X1 g51030(.A (n_5004), .B (n_5014), .C (n_5003), .D (n_5015), .Q
       (n_5791));
  OR4X1 g51031(.A (n_5010), .B (n_5011), .C (n_5012), .D (n_5013), .Q
       (n_5790));
  NA2X1 g51032(.A (n_5408), .B (n_5409), .Q (n_5789));
  NA2X1 g51033(.A (n_5406), .B (n_5407), .Q (n_5788));
  OR4X1 g51034(.A (n_4999), .B (n_5001), .C (n_5000), .D (n_5002), .Q
       (n_5787));
  NA2X1 g51035(.A (n_5404), .B (n_5405), .Q (n_5786));
  NA2X1 g51036(.A (n_5402), .B (n_5403), .Q (n_5785));
  OR4X1 g51037(.A (n_4975), .B (n_4977), .C (n_4976), .D (n_4978), .Q
       (n_5784));
  OR4X1 g51039(.A (n_4915), .B (n_4917), .C (n_4916), .D (n_4914), .Q
       (n_5782));
  OR4X1 g51040(.A (n_4858), .B (n_4859), .C (n_4796), .D (n_4909), .Q
       (n_5781));
  OR4X1 g51044(.A (n_5038), .B (n_4972), .C (n_4986), .D (n_4987), .Q
       (n_5777));
  OR4X1 g51045(.A (n_4970), .B (n_4984), .C (n_4971), .D (n_4985), .Q
       (n_5776));
  OR4X1 g51047(.A (n_4967), .B (n_4968), .C (n_4981), .D (n_4980), .Q
       (n_5774));
  NA2X1 g51048(.A (n_5388), .B (n_5392), .Q (n_5773));
  NA2X1 g51049(.A (n_5387), .B (n_5391), .Q (n_5772));
  OR4X2 g51050(.A (n_4947), .B (n_4946), .C (n_4948), .D (n_4949), .Q
       (n_5771));
  OR4X1 g51051(.A (n_4940), .B (n_4941), .C (n_4942), .D (n_4943), .Q
       (n_5770));
  OR4X1 g51053(.A (n_4930), .B (n_4931), .C (n_4962), .D (n_4963), .Q
       (n_5768));
  OR4X1 g51054(.A (n_4928), .B (n_4929), .C (n_4960), .D (n_4961), .Q
       (n_5767));
  OR4X1 g51055(.A (n_4926), .B (n_4927), .C (n_4958), .D (n_4959), .Q
       (n_5766));
  OR4X1 g51056(.A (n_4924), .B (n_4925), .C (n_4956), .D (n_4957), .Q
       (n_5765));
  OR4X1 g51057(.A (n_4922), .B (n_4923), .C (n_4954), .D (n_4955), .Q
       (n_5764));
  OR4X2 g51060(.A (n_4921), .B (n_4911), .C (n_4953), .D (n_4944), .Q
       (n_5761));
  NA2X1 g51065(.A (n_8473), .B (n_5366), .Q (n_5756));
  NA2X1 g51067(.A (n_5343), .B (n_5345), .Q (n_5754));
  NA2X1 g51073(.A (n_5329), .B (n_5339), .Q (n_5748));
  NA2X1 g51074(.A (n_5328), .B (n_5338), .Q (n_5747));
  NA2X2 g51076(.A (n_5334), .B (n_5335), .Q (n_5745));
  NA2X1 g51077(.A (n_5332), .B (n_5333), .Q (n_5744));
  NA2X1 g51080(.A (n_5324), .B (n_5325), .Q (n_5741));
  NA2X1 g51082(.A (n_5418), .B (instruction[23]), .Q (n_5739));
  NA2X2 g51083(.A (n_5418), .B (instruction[24]), .Q (n_5738));
  NA2X2 g51084(.A (n_5418), .B (instruction[22]), .Q (n_5737));
  NA2X2 g51085(.A (n_5418), .B (n_2431), .Q (n_5736));
  AN22X1 g51086(.A (n_4893), .B (n_7193), .C (n_4891), .D (n_7189), .Q
       (n_5735));
  AN22X1 g51087(.A (n_4893), .B (n_6418), .C (n_4891), .D (n_6414), .Q
       (n_5734));
  AN22X1 g51088(.A (n_4893), .B (n_7224), .C (n_4891), .D (n_7220), .Q
       (n_5733));
  AO22X1 g51090(.A (n_4873), .B (n_6809), .C (n_4882), .D (n_6810), .Q
       (n_5731));
  AN22X1 g51091(.A (n_4500), .B (n_6375), .C (n_4883), .D (n_6376), .Q
       (n_5730));
  AO22X2 g51092(.A (n_4873), .B (n_6995), .C (n_4882), .D (n_6996), .Q
       (n_5729));
  AO22X1 g51093(.A (n_4873), .B (n_6902), .C (n_4882), .D (n_6903), .Q
       (n_5728));
  AN22X1 g51094(.A (n_4901), .B (n_7208), .C (n_4899), .D (n_7204), .Q
       (n_5727));
  AN22X1 g51095(.A (n_4901), .B (n_6433), .C (n_4899), .D (n_6429), .Q
       (n_5726));
  AN22X1 g51096(.A (n_4901), .B (n_7239), .C (n_4899), .D (n_7235), .Q
       (n_5725));
  AN22X1 g51097(.A (n_4901), .B (n_6960), .C (n_4899), .D (n_6956), .Q
       (n_5724));
  AO22X1 g51098(.A (n_4901), .B (n_6805), .C (n_4899), .D (n_6801), .Q
       (n_5723));
  AN22X1 g51100(.A (n_4901), .B (n_6991), .C (n_4899), .D (n_6987), .Q
       (n_5721));
  AO22X1 g51101(.A (n_4901), .B (n_6898), .C (n_4899), .D (n_6894), .Q
       (n_5720));
  AN22X1 g51102(.A (n_4895), .B (n_7209), .C (n_4897), .D (n_7205), .Q
       (n_5719));
  AN22X1 g51103(.A (n_4895), .B (n_6434), .C (n_4897), .D (n_6430), .Q
       (n_5718));
  AN22X1 g51104(.A (n_4895), .B (n_7240), .C (n_4897), .D (n_7236), .Q
       (n_5717));
  AN22X1 g51105(.A (n_4895), .B (n_6961), .C (n_4897), .D (n_6957), .Q
       (n_5716));
  NA2X1 g51106(.A (n_8479), .B (n_8676), .Q (n_5715));
  AO22X1 g51107(.A (n_4895), .B (n_6806), .C (n_4897), .D (n_6802), .Q
       (n_5714));
  NA2X1 g51108(.A (n_5315), .B (n_5314), .Q (n_5713));
  AO22X1 g51110(.A (n_4895), .B (n_6899), .C (n_4897), .D (n_6895), .Q
       (n_5711));
  AO22X1 g51111(.A (n_4878), .B (n_7200), .C (n_4506), .D (n_7201), .Q
       (n_5710));
  AN22X1 g51112(.A (n_4878), .B (n_6425), .C (n_4506), .D (n_6426), .Q
       (n_5709));
  AN22X1 g51113(.A (n_4878), .B (n_7231), .C (n_4506), .D (n_7232), .Q
       (n_5708));
  AO22X1 g51114(.A (n_4878), .B (n_6952), .C (n_4506), .D (n_6953), .Q
       (n_5707));
  AN22X1 g51115(.A (n_4452), .B (n_7212), .C (n_4882), .D (n_7213), .Q
       (n_5706));
  AN22X1 g51116(.A (n_4452), .B (n_6437), .C (n_4882), .D (n_6438), .Q
       (n_5705));
  AN22X1 g51117(.A (n_4452), .B (n_7243), .C (n_4882), .D (n_7244), .Q
       (n_5704));
  ON22X1 g51119(.A (n_4904), .B (n_4564), .C (n_4457), .D (n_4566), .Q
       (n_5702));
  AN22X1 g51123(.A (n_4508), .B (n_7216), .C (n_4502), .D (n_7217), .Q
       (n_5698));
  AN22X1 g51124(.A (n_4508), .B (n_6441), .C (n_4502), .D (n_6442), .Q
       (n_5697));
  AN22X1 g51125(.A (n_4508), .B (n_7247), .C (n_4502), .D (n_7248), .Q
       (n_5696));
  AN22X1 g51126(.A (n_4508), .B (n_6968), .C (n_4502), .D (n_6969), .Q
       (n_5695));
  AN22X1 g51127(.A (n_4901), .B (n_6309), .C (n_4899), .D (n_6305), .Q
       (n_5694));
  NA2X1 g51128(.A (n_5305), .B (n_5304), .Q (n_5693));
  AN22X1 g51129(.A (n_4901), .B (n_6557), .C (n_4899), .D (n_6553), .Q
       (n_5692));
  AO22X1 g51131(.A (n_4901), .B (n_6402), .C (n_4899), .D (n_6398), .Q
       (n_5690));
  AO22X1 g51132(.A (n_4893), .B (n_6790), .C (n_4891), .D (n_6786), .Q
       (n_5689));
  AN22X1 g51133(.A (n_4893), .B (n_6356), .C (n_4891), .D (n_6352), .Q
       (n_5688));
  AN22X1 g51135(.A (n_4893), .B (n_6883), .C (n_4891), .D (n_6879), .Q
       (n_5686));
  AO22X1 g51137(.A (n_4903), .B (n_6789), .C (n_4861), .D (n_6785), .Q
       (n_5684));
  AN22X1 g51138(.A (n_4878), .B (n_6797), .C (n_4506), .D (n_6798), .Q
       (n_5683));
  AN22X1 g51140(.A (n_4878), .B (n_6363), .C (n_4506), .D (n_6364), .Q
       (n_5681));
  NA2X1 g51141(.A (n_5312), .B (n_5313), .Q (n_5680));
  AO22X1 g51143(.A (n_4878), .B (n_6983), .C (n_4506), .D (n_6984), .Q
       (n_5678));
  AO22X1 g51144(.A (n_4895), .B (n_6310), .C (n_4897), .D (n_6306), .Q
       (n_5677));
  AO22X1 g51146(.A (n_4895), .B (n_6279), .C (n_4897), .D (n_6275), .Q
       (n_5675));
  AO22X1 g51147(.A (n_4895), .B (n_6558), .C (n_4897), .D (n_6554), .Q
       (n_5674));
  AN22X1 g51149(.A (n_4893), .B (n_6542), .C (n_4891), .D (n_6538), .Q
       (n_5672));
  NA2X1 g51150(.A (n_5297), .B (n_5296), .Q (n_5671));
  AO22X1 g51151(.A (n_4895), .B (n_6403), .C (n_4897), .D (n_6399), .Q
       (n_5670));
  AN22X1 g51152(.A (n_4893), .B (n_7100), .C (n_4891), .D (n_7096), .Q
       (n_5669));
  AO22X1 g51153(.A (n_4893), .B (n_6387), .C (n_4891), .D (n_6383), .Q
       (n_5668));
  AO22X1 g51154(.A (n_4508), .B (n_6813), .C (n_4502), .D (n_6814), .Q
       (n_5667));
  AN22X1 g51155(.A (n_4508), .B (n_6379), .C (n_4502), .D (n_6380), .Q
       (n_5666));
  AN22X1 g51156(.A (n_4508), .B (n_6999), .C (n_4502), .D (n_7000), .Q
       (n_5665));
  NA2X1 g51158(.A (n_5307), .B (n_5308), .Q (n_5663));
  NA2X1 g51159(.A (n_5306), .B (n_5309), .Q (n_5662));
  NA2X1 g51160(.A (n_5300), .B (n_5303), .Q (n_5661));
  NA2X1 g51161(.A (n_5301), .B (n_5302), .Q (n_5660));
  NA2X1 g51162(.A (n_5298), .B (n_5299), .Q (n_5659));
  NA2X1 g51163(.A (n_5287), .B (n_5288), .Q (n_5658));
  NA2X1 g51164(.A (n_5283), .B (n_5284), .Q (n_5657));
  NA2X1 g51165(.A (n_5280), .B (n_5279), .Q (n_5656));
  NA2X1 g51166(.A (n_5275), .B (n_5276), .Q (n_5655));
  AN22X1 g51168(.A (n_4901), .B (n_7084), .C (n_4899), .D (n_7080), .Q
       (n_5653));
  NA2X1 g51169(.A (n_5268), .B (n_5267), .Q (n_5652));
  NA2X1 g51170(.A (n_5264), .B (n_5263), .Q (n_5651));
  NA2X1 g51171(.A (n_5259), .B (n_5260), .Q (n_5650));
  NA2X1 g51172(.A (n_5258), .B (n_5257), .Q (n_5649));
  NA2X1 g51173(.A (n_5254), .B (n_5255), .Q (n_5648));
  NA2X1 g51174(.A (n_5251), .B (n_5252), .Q (n_5647));
  NA2X1 g51175(.A (n_5250), .B (n_5249), .Q (n_5646));
  AN22X1 g51176(.A (n_4895), .B (n_7085), .C (n_4897), .D (n_7081), .Q
       (n_5645));
  NA2X1 g51177(.A (n_5248), .B (n_5247), .Q (n_5644));
  NA2X1 g51179(.A (n_5285), .B (n_5286), .Q (n_5642));
  NA2X1 g51180(.A (n_5281), .B (n_5282), .Q (n_5641));
  NA2X1 g51181(.A (n_5277), .B (n_5278), .Q (n_5640));
  NA2X1 g51182(.A (n_5273), .B (n_5274), .Q (n_5639));
  NA2X1 g51183(.A (n_5271), .B (n_5272), .Q (n_5638));
  NA2X1 g51184(.A (n_5269), .B (n_5270), .Q (n_5637));
  NA2X1 g51186(.A (n_5261), .B (n_5262), .Q (n_5635));
  AN22X1 g51187(.A (n_4866), .B (n_7198), .C (n_4498), .D (n_7199), .Q
       (n_5634));
  AN22X1 g51188(.A (n_4866), .B (n_6423), .C (n_4498), .D (n_6424), .Q
       (n_5633));
  AN22X1 g51189(.A (n_4866), .B (n_7229), .C (n_4498), .D (n_7230), .Q
       (n_5632));
  AN22X1 g51191(.A (n_4878), .B (n_6301), .C (n_4506), .D (n_6302), .Q
       (n_5630));
  AN22X1 g51192(.A (n_4878), .B (n_6270), .C (n_4506), .D (n_6271), .Q
       (n_5629));
  NA2X1 g51194(.A (n_5292), .B (n_5289), .Q (n_5627));
  AN22X1 g51195(.A (n_4878), .B (n_6394), .C (n_4506), .D (n_6395), .Q
       (n_5626));
  AN22X1 g51197(.A (n_4508), .B (n_6317), .C (n_4502), .D (n_6318), .Q
       (n_5624));
  AO22X1 g51198(.A (n_4500), .B (n_6282), .C (n_4882), .D (n_6283), .Q
       (n_5623));
  AN22X1 g51201(.A (n_4508), .B (n_6565), .C (n_4502), .D (n_6566), .Q
       (n_5620));
  AN22X1 g51202(.A (n_4500), .B (n_7119), .C (n_4883), .D (n_7120), .Q
       (n_5619));
  AN22X1 g51203(.A (n_4508), .B (n_7123), .C (n_4502), .D (n_7124), .Q
       (n_5618));
  AN22X1 g51204(.A (n_4500), .B (n_6406), .C (n_4883), .D (n_6407), .Q
       (n_5617));
  AN22X1 g51205(.A (n_4508), .B (n_6410), .C (n_4502), .D (n_6411), .Q
       (n_5616));
  AN22X1 g51206(.A (n_4868), .B (n_7190), .C (n_4870), .D (n_7191), .Q
       (n_5615));
  AN22X1 g51207(.A (n_4868), .B (n_7221), .C (n_4870), .D (n_7222), .Q
       (n_5614));
  AN22X1 g51208(.A (n_4868), .B (n_6415), .C (n_4870), .D (n_6416), .Q
       (n_5613));
  AO22X1 g51209(.A (n_4868), .B (n_6942), .C (n_4870), .D (n_6943), .Q
       (n_5612));
  AN22X1 g51210(.A (n_4878), .B (n_6921), .C (n_4506), .D (n_6922), .Q
       (n_5611));
  AO22X1 g51211(.A (n_4878), .B (n_6859), .C (n_4506), .D (n_6860), .Q
       (n_5610));
  AO22X1 g51212(.A (n_4878), .B (n_6828), .C (n_4506), .D (n_6829), .Q
       (n_5609));
  NO2X1 g51213(.A (n_5039), .B (n_5040), .Q (n_5608));
  NA2X1 g51214(.A (n_5217), .B (n_5216), .Q (n_5607));
  AO22X1 g51215(.A (n_4878), .B (n_7076), .C (n_4506), .D (n_7077), .Q
       (n_5606));
  NA2X1 g51216(.A (n_5215), .B (n_5214), .Q (n_5605));
  AN22X1 g51217(.A (n_4878), .B (n_6332), .C (n_4506), .D (n_6333), .Q
       (n_5604));
  AN22X1 g51218(.A (n_4893), .B (n_6914), .C (n_4891), .D (n_6910), .Q
       (n_5603));
  NA2X1 g51219(.A (n_5256), .B (n_5213), .Q (n_5602));
  AN22X1 g51221(.A (n_4893), .B (n_7131), .C (n_4891), .D (n_7127), .Q
       (n_5600));
  AN22X1 g51222(.A (n_4893), .B (n_7069), .C (n_4891), .D (n_7065), .Q
       (n_5599));
  AN22X1 g51223(.A (n_4893), .B (n_7007), .C (n_4891), .D (n_7003), .Q
       (n_5598));
  AN22X1 g51226(.A (n_4888), .B (n_6421), .C (n_4884), .D (n_6422), .Q
       (n_5595));
  AN22X1 g51227(.A (n_4888), .B (n_7227), .C (n_4884), .D (n_7228), .Q
       (n_5594));
  AN22X1 g51228(.A (n_4888), .B (n_6948), .C (n_4884), .D (n_6949), .Q
       (n_5593));
  AO22X2 g51230(.A (n_4873), .B (n_6871), .C (n_4882), .D (n_6872), .Q
       (n_5591));
  AN22X1 g51236(.A (n_4500), .B (n_7150), .C (n_4883), .D (n_7151), .Q
       (n_5585));
  AN22X1 g51237(.A (n_4508), .B (n_7154), .C (n_4502), .D (n_7155), .Q
       (n_5584));
  AN22X1 g51238(.A (n_4873), .B (n_7088), .C (n_4883), .D (n_7089), .Q
       (n_5583));
  AN22X1 g51239(.A (n_4508), .B (n_7092), .C (n_4503), .D (n_7093), .Q
       (n_5582));
  AO22X1 g51240(.A (n_4452), .B (n_7026), .C (n_4883), .D (n_7027), .Q
       (n_5581));
  AO22X1 g51242(.A (n_4452), .B (n_6344), .C (n_4883), .D (n_6345), .Q
       (n_5579));
  AO22X1 g51243(.A (n_4508), .B (n_6348), .C (n_4502), .D (n_6349), .Q
       (n_5578));
  NA2X1 g51245(.A (n_5294), .B (n_5295), .Q (n_5576));
  AO22X2 g51246(.A (n_4888), .B (n_6793), .C (n_4884), .D (n_6794), .Q
       (n_5575));
  AN22X1 g51247(.A (n_4888), .B (n_6359), .C (n_4884), .D (n_6360), .Q
       (n_5574));
  AN22X1 g51248(.A (n_4888), .B (n_6979), .C (n_4884), .D (n_6980), .Q
       (n_5573));
  AN22X1 g51249(.A (n_4866), .B (n_6547), .C (n_4498), .D (n_6548), .Q
       (n_5572));
  AN22X1 g51250(.A (n_4866), .B (n_6795), .C (n_4498), .D (n_6796), .Q
       (n_5571));
  AN22X1 g51251(.A (n_4866), .B (n_6392), .C (n_4498), .D (n_6393), .Q
       (n_5570));
  AO22X1 g51252(.A (n_4866), .B (n_6361), .C (n_4498), .D (n_6362), .Q
       (n_5569));
  AN22X1 g51254(.A (n_4866), .B (n_6888), .C (n_4498), .D (n_6889), .Q
       (n_5567));
  AN22X1 g51255(.A (n_4868), .B (n_6539), .C (n_4870), .D (n_6540), .Q
       (n_5566));
  AN22X1 g51256(.A (n_4868), .B (n_6787), .C (n_4870), .D (n_6788), .Q
       (n_5565));
  AN22X1 g51257(.A (n_4868), .B (n_6384), .C (n_4870), .D (n_6385), .Q
       (n_5564));
  AO22X1 g51258(.A (n_4868), .B (n_6353), .C (n_4870), .D (n_6354), .Q
       (n_5563));
  AO22X1 g51259(.A (n_4868), .B (n_6973), .C (n_4870), .D (n_6974), .Q
       (n_5562));
  AN22X1 g51260(.A (n_4868), .B (n_6880), .C (n_4870), .D (n_6881), .Q
       (n_5561));
  AN22X1 g51261(.A (n_4866), .B (n_6299), .C (n_4498), .D (n_6300), .Q
       (n_5560));
  AO22X1 g51262(.A (n_4866), .B (n_6826), .C (n_4497), .D (n_6827), .Q
       (n_5559));
  AN22X1 g51263(.A (n_4866), .B (n_6268), .C (n_4498), .D (n_6269), .Q
       (n_5558));
  AO22X1 g51264(.A (n_4866), .B (n_7136), .C (n_4497), .D (n_7137), .Q
       (n_5557));
  AN22X1 g51265(.A (n_4866), .B (n_7105), .C (n_4498), .D (n_7106), .Q
       (n_5556));
  AO22X1 g51266(.A (n_4866), .B (n_6330), .C (n_4497), .D (n_6331), .Q
       (n_5555));
  AO22X1 g51267(.A (n_4866), .B (n_6919), .C (n_4497), .D (n_6920), .Q
       (n_5554));
  NA2X1 g51268(.A (n_5243), .B (n_5244), .Q (n_5553));
  AN22X1 g51269(.A (n_4868), .B (n_6260), .C (n_4870), .D (n_6261), .Q
       (n_5552));
  AO22X1 g51270(.A (n_4868), .B (n_7128), .C (n_4870), .D (n_7129), .Q
       (n_5551));
  AN22X1 g51271(.A (n_4868), .B (n_7097), .C (n_4870), .D (n_7098), .Q
       (n_5550));
  AO22X1 g51272(.A (n_4868), .B (n_6322), .C (n_4870), .D (n_6323), .Q
       (n_5549));
  NA2X1 g51273(.A (n_5241), .B (n_5242), .Q (n_5548));
  AN22X1 g51274(.A (n_4868), .B (n_6291), .C (n_4870), .D (n_6292), .Q
       (n_5547));
  NA2X1 g51275(.A (n_5225), .B (n_5224), .Q (n_5546));
  NA2X1 g51276(.A (n_5223), .B (n_5222), .Q (n_5545));
  NA2X1 g51277(.A (n_5221), .B (n_5220), .Q (n_5544));
  AO22X2 g51279(.A (n_4888), .B (n_6390), .C (n_4884), .D (n_6391), .Q
       (n_5542));
  AN22X1 g51280(.A (n_4893), .B (n_7162), .C (n_4891), .D (n_7158), .Q
       (n_5541));
  ON22X1 g51281(.A (n_4902), .B (n_4547), .C (n_4900), .D (n_4549), .Q
       (n_5540));
  NO2X1 g51282(.A (n_5195), .B (n_5196), .Q (n_5539));
  NO2X1 g51283(.A (n_5191), .B (n_5192), .Q (n_5538));
  ON22X1 g51285(.A (n_4896), .B (n_4551), .C (n_4898), .D (n_4541), .Q
       (n_5536));
  OA22X1 g51286(.A (n_4896), .B (n_4550), .C (n_4898), .D (n_4552), .Q
       (n_5535));
  ON22X1 g51287(.A (n_4904), .B (n_4548), .C (n_4457), .D (n_4538), .Q
       (n_5534));
  NA2X1 g51288(.A (n_5201), .B (n_5202), .Q (n_5533));
  AN22X1 g51289(.A (n_4888), .B (n_6917), .C (n_4884), .D (n_6918), .Q
       (n_5532));
  AN22X1 g51290(.A (n_4888), .B (n_6855), .C (n_4884), .D (n_6856), .Q
       (n_5531));
  AN22X1 g51291(.A (n_4888), .B (n_6824), .C (n_4884), .D (n_6825), .Q
       (n_5530));
  NO2X1 g51292(.A (n_5193), .B (n_5194), .Q (n_5529));
  AN22X1 g51293(.A (n_4888), .B (n_7165), .C (n_4884), .D (n_7166), .Q
       (n_5528));
  NA2X1 g51294(.A (n_5211), .B (n_5210), .Q (n_5527));
  NA2X1 g51295(.A (n_5209), .B (n_5208), .Q (n_5526));
  NA2X1 g51297(.A (n_5207), .B (n_5206), .Q (n_5524));
  NA2X1 g51298(.A (n_5205), .B (n_5204), .Q (n_5523));
  AO22X2 g51299(.A (n_4868), .B (n_7066), .C (n_4870), .D (n_7067), .Q
       (n_5522));
  AO22X1 g51300(.A (n_4868), .B (n_7004), .C (n_4870), .D (n_7005), .Q
       (n_5521));
  NO2X1 g51301(.A (n_5187), .B (n_5175), .Q (n_5520));
  NO2X1 g51302(.A (n_5178), .B (n_5184), .Q (n_5519));
  NO2X1 g51303(.A (n_5186), .B (n_5173), .Q (n_5518));
  NO2X1 g51305(.A (n_5185), .B (n_5171), .Q (n_5516));
  AN22X1 g51307(.A (n_4893), .B (n_6759), .C (n_4891), .D (n_6755), .Q
       (n_5514));
  NO2X1 g51308(.A (n_5174), .B (n_5181), .Q (n_5513));
  AN22X1 g51309(.A (n_4893), .B (n_6728), .C (n_4891), .D (n_6724), .Q
       (n_5512));
  NA2X1 g51310(.A (n_5172), .B (n_5180), .Q (n_5511));
  AN22X1 g51311(.A (n_4893), .B (n_6697), .C (n_4891), .D (n_6693), .Q
       (n_5510));
  NA2X1 g51312(.A (n_5170), .B (n_5179), .Q (n_5509));
  NA2X1 g51313(.A (n_5168), .B (n_5169), .Q (n_5508));
  AN22X1 g51314(.A (n_4893), .B (n_7038), .C (n_4891), .D (n_7034), .Q
       (n_5507));
  AN22X1 g51316(.A (n_4878), .B (n_7045), .C (n_4506), .D (n_7046), .Q
       (n_5505));
  AN22X1 g51317(.A (n_4878), .B (n_6735), .C (n_4506), .D (n_6736), .Q
       (n_5504));
  AN22X1 g51318(.A (n_4878), .B (n_6704), .C (n_4506), .D (n_6705), .Q
       (n_5503));
  AN22X1 g51319(.A (n_4878), .B (n_6673), .C (n_4506), .D (n_6674), .Q
       (n_5502));
  ON22X1 g51320(.A (n_4887), .B (n_4543), .C (n_4885), .D (n_4542), .Q
       (n_5501));
  AN22X1 g51321(.A (n_4888), .B (n_7041), .C (n_4884), .D (n_7042), .Q
       (n_5500));
  AO22X1 g51326(.A (n_4508), .B (n_6720), .C (n_4876), .D (n_6721), .Q
       (n_5495));
  AO22X1 g51327(.A (n_4508), .B (n_6689), .C (n_4502), .D (n_6690), .Q
       (n_5494));
  NA2X4 g51328(.A (n_4462), .B (n_4712), .Q (n_7692));
  NO2X1 g51329(.A (n_5166), .B (n_5167), .Q (n_5493));
  NA2X1 g51330(.A (n_5164), .B (n_5165), .Q (n_5492));
  AO22X2 g51331(.A (n_4866), .B (n_7074), .C (n_4498), .D (n_7075), .Q
       (n_5491));
  AO22X1 g51332(.A (n_4866), .B (n_7012), .C (n_4497), .D (n_7013), .Q
       (n_5490));
  AN22X1 g51333(.A (n_4886), .B (n_6731), .C (n_4884), .D (n_6732), .Q
       (n_5489));
  AN22X1 g51334(.A (n_4888), .B (n_6700), .C (n_4884), .D (n_6701), .Q
       (n_5488));
  AO22X1 g51335(.A (n_4886), .B (n_6669), .C (n_4884), .D (n_6670), .Q
       (n_5487));
  NA2X1 g51336(.A (n_5148), .B (n_5147), .Q (n_5486));
  NA2X1 g51337(.A (n_5146), .B (n_5145), .Q (n_5485));
  ON22X1 g51338(.A (n_4869), .B (n_4540), .C (n_4871), .D (n_4539), .Q
       (n_5484));
  NA2X1 g51339(.A (n_5162), .B (n_5163), .Q (n_5483));
  NA2X1 g51340(.A (n_5153), .B (n_5143), .Q (n_5482));
  NA2X1 g51341(.A (n_5152), .B (n_5150), .Q (n_5481));
  NA2X1 g51342(.A (n_5151), .B (n_5149), .Q (n_5480));
  NO2X1 g51344(.A (n_5134), .B (n_5135), .Q (n_5478));
  NA2X1 g51345(.A (n_5132), .B (n_5133), .Q (n_5477));
  NA2X1 g51346(.A (n_5130), .B (n_5131), .Q (n_5476));
  NA2X1 g51347(.A (n_5126), .B (n_5129), .Q (n_5475));
  NO2X1 g51348(.A (n_5140), .B (n_5141), .Q (n_5474));
  NA2X1 g51350(.A (n_5136), .B (n_5137), .Q (n_5472));
  NA2X1 g51353(.A (n_5124), .B (n_5127), .Q (n_5469));
  NA2X1 g51354(.A (n_5125), .B (n_5128), .Q (n_5468));
  NO2X1 g51356(.A (n_5122), .B (n_5093), .Q (n_5466));
  AN22X1 g51357(.A (n_4888), .B (n_6576), .C (n_4884), .D (n_6577), .Q
       (n_5465));
  NO2X1 g51358(.A (n_5115), .B (n_5116), .Q (n_5464));
  NO2X1 g51359(.A (n_5113), .B (n_5114), .Q (n_5463));
  OA22X1 g51360(.A (n_4863), .B (n_4545), .C (n_4862), .D (n_4535), .Q
       (n_5462));
  OA22X1 g51361(.A (n_4863), .B (n_4556), .C (n_4862), .D (n_4559), .Q
       (n_5461));
  NO2X1 g51362(.A (n_5092), .B (n_5227), .Q (n_5460));
  NO2X1 g51363(.A (n_5109), .B (n_5110), .Q (n_5459));
  ON22X1 g51364(.A (n_4902), .B (n_4534), .C (n_4900), .D (n_4533), .Q
       (n_5458));
  ON22X1 g51366(.A (n_4902), .B (n_4554), .C (n_4900), .D (n_4560), .Q
       (n_5456));
  ON22X1 g51368(.A (n_4902), .B (n_4555), .C (n_4900), .D (n_4553), .Q
       (n_5454));
  NA2X1 g51369(.A (n_5111), .B (n_5105), .Q (n_5453));
  NO2X2 g51370(.A (n_5103), .B (n_5104), .Q (n_5452));
  ON22X1 g51371(.A (n_4902), .B (n_4529), .C (n_4900), .D (n_4530), .Q
       (n_5451));
  NO2X1 g51372(.A (n_5099), .B (n_5100), .Q (n_5450));
  NO2X1 g51373(.A (n_5096), .B (n_5097), .Q (n_5449));
  NO2X1 g51375(.A (n_5088), .B (n_5089), .Q (n_5447));
  NO2X1 g51376(.A (n_5101), .B (n_5094), .Q (n_5446));
  NO2X1 g51377(.A (n_5095), .B (n_5048), .Q (n_5445));
  NO2X1 g51378(.A (n_5087), .B (n_5047), .Q (n_5444));
  NA2X1 g51379(.A (n_5076), .B (n_5083), .Q (n_5443));
  NO2X1 g51380(.A (n_5075), .B (n_5082), .Q (n_5442));
  NO2X1 g51382(.A (n_5073), .B (n_5080), .Q (n_5440));
  NO2X1 g51384(.A (n_5071), .B (n_5078), .Q (n_5438));
  NA2X1 g51387(.A (n_5068), .B (n_5085), .Q (n_5435));
  NO2X1 g51388(.A (n_5067), .B (n_5084), .Q (n_5434));
  NO2X1 g51390(.A (n_5054), .B (n_5061), .Q (n_5432));
  NO2X2 g51391(.A (n_5053), .B (n_5066), .Q (n_5431));
  NA2X2 g51392(.A (n_5060), .B (n_5051), .Q (n_5430));
  NO2X1 g51395(.A (n_5055), .B (n_5062), .Q (n_5427));
  AN22X1 g51396(.A (n_4889), .B (n_6514), .C (n_4884), .D (n_6515), .Q
       (n_5426));
  NA2X1 g51398(.A (n_5050), .B (n_5058), .Q (n_5424));
  AN22X1 g51399(.A (n_4499), .B (n_6609), .C (n_4497), .D (n_6610), .Q
       (n_5423));
  NO2X1 g51400(.A (n_5041), .B (n_5042), .Q (n_5422));
  NO2X1 g51401(.A (n_5112), .B (n_5046), .Q (n_5421));
  AN22X1 g51403(.A (n_4878), .B (n_7169), .C (n_4506), .D (n_7170), .Q
       (n_5419));
  AN22X1 g51404(.A (n_4484), .B (n_6625), .C (n_4744), .D (n_6626), .Q
       (n_5417));
  AN22X1 g51405(.A (n_4489), .B (n_6435), .C (n_4738), .D (n_6436), .Q
       (n_5416));
  AN22X1 g51408(.A (n_4745), .B (n_6431), .C (n_4488), .D (n_6432), .Q
       (n_5413));
  AN22X1 g51409(.A (n_4484), .B (n_6439), .C (n_4744), .D (n_6440), .Q
       (n_5412));
  ON22X1 g51411(.A (n_4742), .B (n_4565), .C (n_4743), .D (n_4563), .Q
       (n_5410));
  AN21X1 g51412(.A (n_4481), .B (n_6365), .C (n_5009), .Q (n_5409));
  AN22X1 g51413(.A (n_4489), .B (n_6373), .C (n_4738), .D (n_6374), .Q
       (n_5408));
  AN21X1 g51414(.A (n_4481), .B (n_6985), .C (n_5008), .Q (n_5407));
  AN21X1 g51415(.A (n_4489), .B (n_6993), .C (n_5007), .Q (n_5406));
  AN22X1 g51416(.A (n_4745), .B (n_6369), .C (n_4488), .D (n_6370), .Q
       (n_5405));
  AN22X1 g51417(.A (n_4484), .B (n_6377), .C (n_4744), .D (n_6378), .Q
       (n_5404));
  AN22X1 g51418(.A (n_4745), .B (n_6989), .C (n_4488), .D (n_6990), .Q
       (n_5403));
  AN22X1 g51419(.A (n_4484), .B (n_6997), .C (n_4744), .D (n_6998), .Q
       (n_5402));
  AN22X1 g51420(.A (n_4478), .B (n_7194), .C (n_4492), .D (n_7195), .Q
       (n_5401));
  AN22X1 g51421(.A (n_4478), .B (n_7225), .C (n_4492), .D (n_7226), .Q
       (n_5400));
  AN22X1 g51422(.A (n_4478), .B (n_6419), .C (n_4492), .D (n_6420), .Q
       (n_5399));
  AN22X1 g51423(.A (n_4720), .B (n_6357), .C (n_4492), .D (n_6358), .Q
       (n_5398));
  AN22X1 g51424(.A (n_4720), .B (n_6977), .C (n_4492), .D (n_6978), .Q
       (n_5397));
  AN22X1 g51425(.A (n_4478), .B (n_6946), .C (n_4492), .D (n_6947), .Q
       (n_5396));
  AN22X1 g51426(.A (n_4720), .B (n_6884), .C (n_4756), .D (n_6885), .Q
       (n_5395));
  NO2X1 g51427(.A (n_4989), .B (n_4990), .Q (n_5394));
  AN21X1 g51428(.A (n_4489), .B (n_6280), .C (n_4988), .Q (n_5393));
  AN21X1 g51429(.A (n_4481), .B (n_6396), .C (n_4979), .Q (n_5392));
  AN22X1 g51430(.A (n_4489), .B (n_6404), .C (n_4738), .D (n_6405), .Q
       (n_5391));
  AN21X1 g51431(.A (n_4745), .B (n_6276), .C (n_4974), .Q (n_5390));
  AN22X1 g51432(.A (n_4484), .B (n_6284), .C (n_4744), .D (n_6285), .Q
       (n_5389));
  AN22X1 g51433(.A (n_4745), .B (n_6400), .C (n_4488), .D (n_6401), .Q
       (n_5388));
  AN22X1 g51434(.A (n_4484), .B (n_6408), .C (n_4744), .D (n_6409), .Q
       (n_5387));
  OR2X2 g51438(.A (n_4918), .B (n_4919), .Q (n_5383));
  AN22X1 g51439(.A (n_4720), .B (n_6295), .C (n_4492), .D (n_6296), .Q
       (n_5382));
  AN22X1 g51440(.A (n_4720), .B (n_6264), .C (n_4756), .D (n_6265), .Q
       (n_5381));
  AN22X1 g51441(.A (n_4720), .B (n_6791), .C (n_4756), .D (n_6792), .Q
       (n_5380));
  AN22X1 g51442(.A (n_4478), .B (n_6543), .C (n_4756), .D (n_6544), .Q
       (n_5379));
  AN22X1 g51443(.A (n_4720), .B (n_6388), .C (n_4756), .D (n_6389), .Q
       (n_5378));
  AN22X1 g51444(.A (n_4478), .B (n_6853), .C (n_4756), .D (n_6854), .Q
       (n_5377));
  NO2X1 g51445(.A (n_4825), .B (n_4826), .Q (n_5376));
  AN22X1 g51446(.A (n_4478), .B (n_7132), .C (n_4756), .D (n_7133), .Q
       (n_5375));
  AN22X1 g51447(.A (n_4720), .B (n_7101), .C (n_4492), .D (n_7102), .Q
       (n_5374));
  AN22X1 g51448(.A (n_4478), .B (n_6326), .C (n_4756), .D (n_6327), .Q
       (n_5373));
  NO2X1 g51449(.A (n_4833), .B (n_4834), .Q (n_5372));
  NO2X1 g51450(.A (n_4829), .B (n_4830), .Q (n_5371));
  NO2X1 g51453(.A (n_4819), .B (n_4820), .Q (n_5368));
  AN22X1 g51454(.A (n_4478), .B (n_7008), .C (n_4492), .D (n_7009), .Q
       (n_5367));
  NO2X2 g51455(.A (n_4804), .B (n_4805), .Q (n_5366));
  NO2X1 g51459(.A (n_4797), .B (n_4798), .Q (n_5362));
  NO2X1 g51462(.A (n_4839), .B (n_4840), .Q (n_5359));
  OA22X1 g51463(.A (n_4750), .B (n_4546), .C (n_4459), .D (n_4537), .Q
       (n_5358));
  NO2X1 g51464(.A (n_4837), .B (n_4838), .Q (n_5357));
  NO2X1 g51467(.A (n_4813), .B (n_4814), .Q (n_5354));
  NO2X1 g51468(.A (n_4807), .B (n_4812), .Q (n_5353));
  NO2X1 g51469(.A (n_4810), .B (n_4811), .Q (n_5352));
  NO2X1 g51470(.A (n_4808), .B (n_4809), .Q (n_5351));
  OA22X1 g51471(.A (n_4718), .B (n_4544), .C (n_4494), .D (n_4536), .Q
       (n_5350));
  NO2X1 g51472(.A (n_4793), .B (n_4794), .Q (n_5349));
  AN22X1 g51474(.A (n_4478), .B (n_6698), .C (n_4492), .D (n_6699), .Q
       (n_5347));
  AN22X1 g51475(.A (n_4478), .B (n_6667), .C (n_4492), .D (n_6668), .Q
       (n_5346));
  AO21X1 g51476(.A (n_4696), .B (n_8484), .C (n_4907), .Q (n_7671));
  NO2X1 g51477(.A (n_4783), .B (n_4784), .Q (n_5345));
  NO2X1 g51479(.A (n_4786), .B (n_4785), .Q (n_5343));
  AN22X1 g51480(.A (n_4484), .B (n_6594), .C (n_4744), .D (n_6595), .Q
       (n_5342));
  NA2I1X1 g51481(.B (n_4906), .AN (n_4732), .Q (n_7672));
  NA2I1X1 g51482(.B (n_4906), .AN (n_4737), .Q (n_7673));
  NA2I1X1 g51483(.B (n_4906), .AN (n_4736), .Q (n_7674));
  AN22X1 g51484(.A (n_4478), .B (n_6574), .C (n_4492), .D (n_6575), .Q
       (n_5341));
  AO22X1 g51485(.A (n_4478), .B (n_6450), .C (n_4492), .D (n_6451), .Q
       (n_5340));
  NA2X1 g51486(.A (n_4906), .B (n_4734), .Q (n_7677));
  NA2X1 g51487(.A (n_4906), .B (n_4735), .Q (n_7676));
  NA2X1 g51488(.A (n_4906), .B (n_4733), .Q (n_7675));
  AN22X1 g51489(.A (n_4739), .B (n_6644), .C (n_4491), .D (n_6645), .Q
       (n_5339));
  AN22X1 g51490(.A (n_4489), .B (n_6652), .C (n_4738), .D (n_6653), .Q
       (n_5338));
  OA22X2 g51491(.A (n_4740), .B (n_4557), .C (n_4460), .D (n_4558), .Q
       (n_5337));
  AN22X1 g51492(.A (n_4748), .B (n_6621), .C (n_4738), .D (n_6622), .Q
       (n_5336));
  OA22X2 g51493(.A (n_4740), .B (n_4561), .C (n_4460), .D (n_4562), .Q
       (n_5335));
  AN22X1 g51494(.A (n_4489), .B (n_6528), .C (n_4738), .D (n_6529), .Q
       (n_5334));
  AN22X1 g51495(.A (n_4739), .B (n_6489), .C (n_4491), .D (n_6490), .Q
       (n_5333));
  AN22X1 g51496(.A (n_4748), .B (n_6497), .C (n_4738), .D (n_6498), .Q
       (n_5332));
  OA22X2 g51497(.A (n_4480), .B (n_4531), .C (n_4460), .D (n_4532), .Q
       (n_5331));
  AN22X1 g51498(.A (n_4748), .B (n_6466), .C (n_4738), .D (n_6467), .Q
       (n_5330));
  AN22X1 g51499(.A (n_4745), .B (n_6648), .C (n_4488), .D (n_6649), .Q
       (n_5329));
  AN22X1 g51500(.A (n_4484), .B (n_6656), .C (n_4744), .D (n_6657), .Q
       (n_5328));
  AN22X1 g51502(.A (n_4481), .B (n_6427), .C (n_4491), .D (n_6428), .Q
       (n_5326));
  NO2X1 g51503(.A (n_4769), .B (n_4775), .Q (n_5325));
  AN22X1 g51504(.A (n_4484), .B (n_6532), .C (n_4744), .D (n_6533), .Q
       (n_5324));
  NO2X1 g51507(.A (n_4768), .B (n_4776), .Q (n_5321));
  AN22X1 g51508(.A (n_4484), .B (n_6470), .C (n_4744), .D (n_6471), .Q
       (n_5320));
  AO21X1 g51511(.A (n_4696), .B (instruction[22]), .C (n_4907), .Q
       (n_7669));
  AO21X1 g51512(.A (n_4696), .B (instruction[23]), .C (n_4907), .Q
       (n_7678));
  NA2X1 g51515(.A (n_4897), .B (n_6368), .Q (n_5315));
  NA2X1 g51516(.A (n_4895), .B (n_6372), .Q (n_5314));
  NA2X1 g51517(.A (n_4861), .B (n_6971), .Q (n_5313));
  NA2X1 g51518(.A (n_4903), .B (n_6975), .Q (n_5312));
  NA2X1 g51521(.A (n_4861), .B (n_6537), .Q (n_5309));
  NA2X1 g51522(.A (n_4861), .B (n_6258), .Q (n_5308));
  NA2X1 g51523(.A (n_4903), .B (n_6262), .Q (n_5307));
  NA2X1 g51524(.A (n_4903), .B (n_6541), .Q (n_5306));
  NA2X1 g51525(.A (n_4899), .B (n_6274), .Q (n_5305));
  NA2X1 g51526(.A (n_4901), .B (n_6278), .Q (n_5304));
  NA2X1 g51527(.A (n_4861), .B (n_6382), .Q (n_5303));
  NA2X1 g51528(.A (n_4861), .B (n_7095), .Q (n_5302));
  NA2X1 g51529(.A (n_4903), .B (n_7099), .Q (n_5301));
  NA2X1 g51530(.A (n_4903), .B (n_6386), .Q (n_5300));
  NA2X1 g51531(.A (n_4861), .B (n_6289), .Q (n_5299));
  NA2X1 g51532(.A (n_4903), .B (n_6293), .Q (n_5298));
  NA2X1 g51533(.A (n_4897), .B (n_7112), .Q (n_5297));
  NA2X1 g51534(.A (n_4895), .B (n_7116), .Q (n_5296));
  NA2X1 g51535(.A (n_4884), .B (n_6887), .Q (n_5295));
  NA2X1 g51536(.A (n_4888), .B (n_6886), .Q (n_5294));
  NA2X1 g51539(.A (n_4506), .B (n_7108), .Q (n_5292));
  NA2X1 g51542(.A (n_4878), .B (n_7107), .Q (n_5289));
  NA2X1 g51543(.A (n_4899), .B (n_6925), .Q (n_5288));
  NA2X1 g51544(.A (n_4901), .B (n_6929), .Q (n_5287));
  NA2X1 g51545(.A (n_4861), .B (n_6847), .Q (n_5286));
  NA2X1 g51546(.A (n_4903), .B (n_6851), .Q (n_5285));
  NA2X1 g51547(.A (n_4899), .B (n_6863), .Q (n_5284));
  NA2X1 g51548(.A (n_4901), .B (n_6867), .Q (n_5283));
  NA2X1 g51549(.A (n_4861), .B (n_6816), .Q (n_5282));
  NA2X1 g51550(.A (n_4903), .B (n_6820), .Q (n_5281));
  NA2X1 g51551(.A (n_4899), .B (n_6832), .Q (n_5280));
  NA2X1 g51552(.A (n_4901), .B (n_6836), .Q (n_5279));
  NA2X1 g51553(.A (n_4861), .B (n_7157), .Q (n_5278));
  NA2X1 g51554(.A (n_4903), .B (n_7161), .Q (n_5277));
  NA2X1 g51555(.A (n_4899), .B (n_7173), .Q (n_5276));
  NA2X1 g51556(.A (n_4901), .B (n_7177), .Q (n_5275));
  NA2X1 g51557(.A (n_4861), .B (n_7126), .Q (n_5274));
  NA2X1 g51558(.A (n_4903), .B (n_7130), .Q (n_5273));
  NA2X1 g51559(.A (n_4861), .B (n_7064), .Q (n_5272));
  NA2X1 g51560(.A (n_4903), .B (n_7068), .Q (n_5271));
  NA2X1 g51561(.A (n_4861), .B (n_7002), .Q (n_5270));
  NA2X1 g51562(.A (n_4903), .B (n_7006), .Q (n_5269));
  NA2X1 g51563(.A (n_4899), .B (n_7018), .Q (n_5268));
  NA2X1 g51564(.A (n_4901), .B (n_7022), .Q (n_5267));
  NA2X1 g51567(.A (n_4899), .B (n_6336), .Q (n_5264));
  NA2X1 g51568(.A (n_4901), .B (n_6340), .Q (n_5263));
  NA2X1 g51569(.A (n_4861), .B (n_6909), .Q (n_5262));
  NA2X1 g51570(.A (n_4903), .B (n_6913), .Q (n_5261));
  NA2X1 g51571(.A (n_4897), .B (n_6926), .Q (n_5260));
  NA2X1 g51572(.A (n_4895), .B (n_6930), .Q (n_5259));
  NA2X1 g51573(.A (n_4897), .B (n_6864), .Q (n_5258));
  NA2X1 g51574(.A (n_4895), .B (n_6868), .Q (n_5257));
  NA2X1 g51575(.A (n_4893), .B (n_6852), .Q (n_5256));
  NA2X1 g51576(.A (n_4897), .B (n_6833), .Q (n_5255));
  NA2X1 g51577(.A (n_4895), .B (n_6837), .Q (n_5254));
  NA2X1 g51579(.A (n_4897), .B (n_7174), .Q (n_5252));
  NA2X1 g51580(.A (n_4895), .B (n_7178), .Q (n_5251));
  NA2X1 g51581(.A (n_4897), .B (n_7143), .Q (n_5250));
  NA2X1 g51582(.A (n_4895), .B (n_7147), .Q (n_5249));
  NA2X1 g51583(.A (n_4897), .B (n_7019), .Q (n_5248));
  NA2X1 g51584(.A (n_4895), .B (n_7023), .Q (n_5247));
  NA2X1 g51587(.A (n_4870), .B (n_6819), .Q (n_5244));
  NA2X1 g51588(.A (n_4868), .B (n_6818), .Q (n_5243));
  NA2X1 g51589(.A (n_4870), .B (n_6912), .Q (n_5242));
  NA2X1 g51590(.A (n_4868), .B (n_6911), .Q (n_5241));
  NA2X4 g51600(.A (n_4908), .B (n_4684), .Q (n_5418));
  INX1 g51601(.A (n_8479), .Q (n_5230));
  INX1 g51602(.A (n_5229), .Q (n_5228));
  NO2I1X1 g51603(.B (n_4869), .AN (n_6477), .Q (n_5227));
  NA2X1 g51605(.A (n_4884), .B (n_6298), .Q (n_5225));
  NA2X1 g51606(.A (n_4888), .B (n_6297), .Q (n_5224));
  NA2X1 g51607(.A (n_4884), .B (n_6267), .Q (n_5223));
  NA2X1 g51608(.A (n_4888), .B (n_6266), .Q (n_5222));
  NA2X1 g51609(.A (n_4884), .B (n_6546), .Q (n_5221));
  NA2X1 g51610(.A (n_4888), .B (n_6545), .Q (n_5220));
  NA2X1 g51613(.A (n_4506), .B (n_7139), .Q (n_5217));
  NA2X1 g51614(.A (n_4878), .B (n_7138), .Q (n_5216));
  NA2X1 g51615(.A (n_4506), .B (n_7015), .Q (n_5215));
  NA2X1 g51616(.A (n_4878), .B (n_7014), .Q (n_5214));
  NA2X1 g51617(.A (n_4891), .B (n_6848), .Q (n_5213));
  AO21X2 g51619(.A (n_4696), .B (n_2431), .C (n_4907), .Q (n_7693));
  NA2X2 g51620(.A (n_4906), .B (n_4711), .Q (n_7670));
  NA2X1 g51621(.A (n_4884), .B (n_7135), .Q (n_5211));
  NA2X1 g51622(.A (n_4888), .B (n_7134), .Q (n_5210));
  NA2X1 g51623(.A (n_4884), .B (n_7073), .Q (n_5209));
  NA2X1 g51624(.A (n_4888), .B (n_7072), .Q (n_5208));
  NA2X1 g51625(.A (n_4884), .B (n_7011), .Q (n_5207));
  NA2X1 g51626(.A (n_4888), .B (n_7010), .Q (n_5206));
  NA2X1 g51627(.A (n_4884), .B (n_6329), .Q (n_5205));
  NA2X1 g51628(.A (n_4888), .B (n_6328), .Q (n_5204));
  NA2X1 g51630(.A (n_4861), .B (n_7033), .Q (n_5202));
  NA2X1 g51631(.A (n_4903), .B (n_7037), .Q (n_5201));
  NO2I1X1 g51632(.B (n_4900), .AN (n_7049), .Q (n_5200));
  NO2I1X1 g51633(.B (n_4902), .AN (n_7053), .Q (n_5199));
  NA2X1 g51634(.A (n_4870), .B (n_6850), .Q (n_5198));
  NA2X1 g51635(.A (n_4868), .B (n_6849), .Q (n_5197));
  NO2I1X1 g51638(.B (n_4507), .AN (n_6779), .Q (n_5196));
  NO2I1X1 g51639(.B (n_4874), .AN (n_6778), .Q (n_5195));
  NO2I1X1 g51640(.B (n_4504), .AN (n_6783), .Q (n_5194));
  NO2I1X1 g51641(.B (n_4463), .AN (n_6782), .Q (n_5193));
  NO2I1X1 g51642(.B (n_4507), .AN (n_7058), .Q (n_5192));
  NO2I1X1 g51643(.B (n_4874), .AN (n_7057), .Q (n_5191));
  NO2I1X1 g51644(.B (n_4504), .AN (n_7062), .Q (n_5190));
  NO2I1X1 g51648(.B (n_4904), .AN (n_6727), .Q (n_5187));
  NO2I1X1 g51649(.B (n_4904), .AN (n_6696), .Q (n_5186));
  NO2I1X1 g51650(.B (n_4904), .AN (n_6665), .Q (n_5185));
  NO2I1X1 g51651(.B (n_4900), .AN (n_6739), .Q (n_5184));
  NA2X1 g51652(.A (n_4899), .B (n_6708), .Q (n_5183));
  NA2X1 g51653(.A (n_4899), .B (n_6677), .Q (n_5182));
  NO2I1X1 g51654(.B (n_4898), .AN (n_6740), .Q (n_5181));
  NA2X1 g51655(.A (n_4897), .B (n_6709), .Q (n_5180));
  NA2X1 g51656(.A (n_4897), .B (n_6678), .Q (n_5179));
  NO2I1X1 g51657(.B (n_4902), .AN (n_6743), .Q (n_5178));
  NA2X1 g51658(.A (n_4901), .B (n_6712), .Q (n_5177));
  NA2X1 g51659(.A (n_4901), .B (n_6681), .Q (n_5176));
  NO2I1X1 g51660(.B (n_4457), .AN (n_6723), .Q (n_5175));
  NO2I1X1 g51661(.B (n_4896), .AN (n_6744), .Q (n_5174));
  NO2I1X1 g51662(.B (n_4457), .AN (n_6692), .Q (n_5173));
  NA2X1 g51663(.A (n_4895), .B (n_6713), .Q (n_5172));
  NO2I1X1 g51664(.B (n_4457), .AN (n_6661), .Q (n_5171));
  NA2X1 g51665(.A (n_4895), .B (n_6682), .Q (n_5170));
  NA2X1 g51666(.A (n_4891), .B (n_6662), .Q (n_5169));
  NA2X1 g51667(.A (n_4893), .B (n_6666), .Q (n_5168));
  NO2I1X1 g51668(.B (n_4862), .AN (n_6858), .Q (n_5167));
  NO2I1X1 g51669(.B (n_4863), .AN (n_6857), .Q (n_5166));
  NA2X1 g51670(.A (n_4498), .B (n_7168), .Q (n_5165));
  NA2X1 g51671(.A (n_4866), .B (n_7167), .Q (n_5164));
  NA2X1 g51672(.A (n_4870), .B (n_7036), .Q (n_5163));
  NA2X1 g51673(.A (n_4868), .B (n_7035), .Q (n_5162));
  NO2I1X1 g51674(.B (n_4881), .AN (n_6748), .Q (n_5161));
  NO2I1X1 g51675(.B (n_4874), .AN (n_6747), .Q (n_5160));
  NO2I1X1 g51676(.B (n_4504), .AN (n_6752), .Q (n_5159));
  NA2X1 g51678(.A (n_4883), .B (n_6717), .Q (n_5157));
  NA2X1 g51679(.A (n_4500), .B (n_6716), .Q (n_5156));
  NA2X1 g51680(.A (n_4883), .B (n_6686), .Q (n_5155));
  NA2X1 g51681(.A (n_4500), .B (n_6685), .Q (n_5154));
  NA2X1 g51682(.A (n_4903), .B (n_6572), .Q (n_5153));
  NA2X1 g51683(.A (n_4899), .B (n_6584), .Q (n_5152));
  NA2X1 g51684(.A (n_4897), .B (n_6585), .Q (n_5151));
  NA2X1 g51685(.A (n_4901), .B (n_6588), .Q (n_5150));
  NA2X1 g51686(.A (n_4895), .B (n_6589), .Q (n_5149));
  NA2X1 g51687(.A (n_4498), .B (n_6765), .Q (n_5148));
  NA2X1 g51688(.A (n_4866), .B (n_6764), .Q (n_5147));
  NA2X1 g51689(.A (n_4498), .B (n_7044), .Q (n_5146));
  NA2X1 g51690(.A (n_4866), .B (n_7043), .Q (n_5145));
  NA2X1 g51692(.A (n_4861), .B (n_6568), .Q (n_5143));
  NO2I1X1 g51694(.B (n_4862), .AN (n_6734), .Q (n_5141));
  NO2I1X1 g51695(.B (n_4863), .AN (n_6733), .Q (n_5140));
  NA2X1 g51698(.A (n_4498), .B (n_6672), .Q (n_5137));
  NA2X1 g51699(.A (n_4866), .B (n_6671), .Q (n_5136));
  NO2I1X1 g51700(.B (n_4871), .AN (n_6726), .Q (n_5135));
  NO2I1X1 g51701(.B (n_4869), .AN (n_6725), .Q (n_5134));
  NA2X1 g51702(.A (n_4870), .B (n_6695), .Q (n_5133));
  NA2X1 g51703(.A (n_4868), .B (n_6694), .Q (n_5132));
  NA2X1 g51704(.A (n_4870), .B (n_6664), .Q (n_5131));
  NA2X1 g51705(.A (n_4868), .B (n_6663), .Q (n_5130));
  NA2X1 g51706(.A (n_4506), .B (n_6581), .Q (n_5129));
  NA2X1 g51707(.A (n_4503), .B (n_6597), .Q (n_5128));
  NA2X1 g51708(.A (n_4883), .B (n_6593), .Q (n_5127));
  NA2X1 g51709(.A (n_4878), .B (n_6580), .Q (n_5126));
  NA2X1 g51710(.A (n_4508), .B (n_6596), .Q (n_5125));
  NA2X1 g51711(.A (n_4452), .B (n_6592), .Q (n_5124));
  NO2I1X1 g51712(.B (n_4892), .AN (n_6631), .Q (n_5123));
  NO2I1X1 g51713(.B (n_4892), .AN (n_6507), .Q (n_5122));
  NO2I1X1 g51714(.B (n_4892), .AN (n_6476), .Q (n_5121));
  NO2I1X1 g51719(.B (n_4871), .AN (n_6633), .Q (n_5116));
  NO2I1X1 g51720(.B (n_4869), .AN (n_6632), .Q (n_5115));
  NO2I1X1 g51721(.B (n_4871), .AN (n_6509), .Q (n_5114));
  NO2I1X1 g51722(.B (n_4869), .AN (n_6508), .Q (n_5113));
  NO2I1X2 g51723(.B (n_4863), .AN (n_6454), .Q (n_5112));
  NA2X1 g51724(.A (n_4899), .B (n_6491), .Q (n_5111));
  NO2I1X1 g51725(.B (n_4457), .AN (n_6630), .Q (n_5110));
  NO2I1X1 g51726(.B (n_4904), .AN (n_6634), .Q (n_5109));
  NO2I1X1 g51727(.B (n_4457), .AN (n_6599), .Q (n_5108));
  NO2I1X1 g51728(.B (n_4904), .AN (n_6603), .Q (n_5107));
  NO2I1X1 g51729(.B (n_4904), .AN (n_6510), .Q (n_5106));
  NA2X1 g51732(.A (n_4901), .B (n_6495), .Q (n_5105));
  NO2I1X1 g51733(.B (n_4457), .AN (n_6444), .Q (n_5104));
  NO2I1X1 g51734(.B (n_4904), .AN (n_6448), .Q (n_5103));
  NO2I1X1 g51735(.B (n_4457), .AN (n_6506), .Q (n_5102));
  NO2I1X1 g51736(.B (n_4896), .AN (n_6527), .Q (n_5101));
  NO2I1X1 g51737(.B (n_4898), .AN (n_6647), .Q (n_5100));
  NO2I1X1 g51738(.B (n_4896), .AN (n_6651), .Q (n_5099));
  NO2I1X1 g51740(.B (n_4898), .AN (n_6616), .Q (n_5097));
  NO2I1X1 g51741(.B (n_4896), .AN (n_6620), .Q (n_5096));
  NO2I1X1 g51742(.B (n_4894), .AN (n_6604), .Q (n_5095));
  NO2I1X1 g51743(.B (n_4898), .AN (n_6523), .Q (n_5094));
  NO2I1X1 g51744(.B (n_4894), .AN (n_6511), .Q (n_5093));
  NO2I1X1 g51745(.B (n_4894), .AN (n_6480), .Q (n_5092));
  NO2I1X1 g51746(.B (n_4898), .AN (n_6492), .Q (n_5091));
  NO2I1X1 g51747(.B (n_4896), .AN (n_6496), .Q (n_5090));
  NO2I1X1 g51748(.B (n_4898), .AN (n_6461), .Q (n_5089));
  NO2I1X1 g51749(.B (n_4896), .AN (n_6465), .Q (n_5088));
  NO2I1X1 g51750(.B (n_4894), .AN (n_6449), .Q (n_5087));
  NO2I1X2 g51751(.B (n_4507), .AN (n_6500), .Q (n_5086));
  NA2X1 g51752(.A (n_4883), .B (n_6469), .Q (n_5085));
  NO2I1X1 g51753(.B (n_4504), .AN (n_6473), .Q (n_5084));
  NA2X1 g51754(.A (n_4883), .B (n_6655), .Q (n_5083));
  NO2I1X1 g51755(.B (n_4504), .AN (n_6659), .Q (n_5082));
  NO2I1X1 g51757(.B (n_4504), .AN (n_6628), .Q (n_5080));
  NA2X1 g51758(.A (n_4883), .B (n_6531), .Q (n_5079));
  NO2I1X1 g51759(.B (n_4504), .AN (n_6535), .Q (n_5078));
  NA2X1 g51761(.A (n_4452), .B (n_6654), .Q (n_5076));
  NO2I1X1 g51762(.B (n_4463), .AN (n_6658), .Q (n_5075));
  NO2I1X1 g51764(.B (n_4463), .AN (n_6627), .Q (n_5073));
  NA2X1 g51765(.A (n_4452), .B (n_6530), .Q (n_5072));
  NO2I1X1 g51766(.B (n_4463), .AN (n_6534), .Q (n_5071));
  NO2I1X2 g51767(.B (n_4874), .AN (n_6499), .Q (n_5070));
  NA2X1 g51769(.A (n_4452), .B (n_6468), .Q (n_5068));
  NO2I1X1 g51770(.B (n_4463), .AN (n_6472), .Q (n_5067));
  NO2I1X2 g51771(.B (n_4505), .AN (n_6519), .Q (n_5066));
  NO2I1X1 g51775(.B (n_4885), .AN (n_6608), .Q (n_5062));
  NO2I1X1 g51776(.B (n_4505), .AN (n_6612), .Q (n_5061));
  NA2X1 g51777(.A (n_4506), .B (n_6488), .Q (n_5060));
  NA2X2 g51779(.A (n_4884), .B (n_6453), .Q (n_5058));
  NO2I1X1 g51782(.B (n_4509), .AN (n_6607), .Q (n_5055));
  NO2I1X1 g51783(.B (n_4879), .AN (n_6611), .Q (n_5054));
  NO2I1X1 g51784(.B (n_4879), .AN (n_6518), .Q (n_5053));
  NA2X1 g51786(.A (n_4878), .B (n_6487), .Q (n_5051));
  NA2X1 g51787(.A (n_4889), .B (n_6452), .Q (n_5050));
  NO2I1X1 g51789(.B (n_4892), .AN (n_6600), .Q (n_5048));
  NO2I1X1 g51790(.B (n_4892), .AN (n_6445), .Q (n_5047));
  NO2I1X1 g51791(.B (n_4862), .AN (n_6455), .Q (n_5046));
  NO2I1X1 g51792(.B (n_4862), .AN (n_6486), .Q (n_5045));
  NO2I1X1 g51793(.B (n_4871), .AN (n_6602), .Q (n_5044));
  NO2I1X1 g51794(.B (n_4869), .AN (n_6601), .Q (n_5043));
  NO2I1X1 g51795(.B (n_4871), .AN (n_6478), .Q (n_5042));
  NO2I1X2 g51796(.B (n_4863), .AN (n_6485), .Q (n_5041));
  NO2I1X1 g51797(.B (n_4871), .AN (n_6447), .Q (n_5040));
  NO2I1X1 g51798(.B (n_4869), .AN (n_6446), .Q (n_5039));
  NO2X2 g51800(.A (n_4905), .B (jal_type), .Q (n_5229));
  NO2I1X1 g51801(.B (n_4485), .AN (n_6555), .Q (n_5038));
  NO2I1X1 g51802(.B (n_4753), .AN (n_7203), .Q (n_5037));
  NO2I1X1 g51803(.B (n_4459), .AN (n_7211), .Q (n_5036));
  NO2I1X1 g51804(.B (n_4750), .AN (n_7210), .Q (n_5035));
  NO2I1X1 g51805(.B (n_4753), .AN (n_7234), .Q (n_5034));
  NO2I1X1 g51808(.B (n_4753), .AN (n_6955), .Q (n_5031));
  NO2I1X1 g51809(.B (n_4482), .AN (n_6954), .Q (n_5030));
  NO2I1X1 g51810(.B (n_4459), .AN (n_6963), .Q (n_5029));
  NO2I1X1 g51811(.B (n_4490), .AN (n_6962), .Q (n_5028));
  NO2I1X1 g51812(.B (n_4747), .AN (n_7207), .Q (n_5027));
  NO2I1X1 g51813(.B (n_4485), .AN (n_7206), .Q (n_5026));
  NO2I1X1 g51814(.B (n_4743), .AN (n_7215), .Q (n_5025));
  NO2I1X1 g51815(.B (n_4742), .AN (n_7214), .Q (n_5024));
  NO2I1X1 g51818(.B (n_4747), .AN (n_6959), .Q (n_5021));
  NO2I1X1 g51819(.B (n_4486), .AN (n_6958), .Q (n_5020));
  NO2I1X1 g51820(.B (n_4743), .AN (n_6967), .Q (n_5019));
  NO2I1X1 g51821(.B (n_4742), .AN (n_6966), .Q (n_5018));
  NO2I1X1 g51822(.B (n_4490), .AN (n_6900), .Q (n_5017));
  NO2I1X1 g51823(.B (n_4459), .AN (n_6901), .Q (n_5016));
  NO2I1X1 g51824(.B (n_4753), .AN (n_6893), .Q (n_5015));
  NO2I1X1 g51825(.B (n_4482), .AN (n_6892), .Q (n_5014));
  NO2I1X1 g51826(.B (n_4753), .AN (n_6800), .Q (n_5013));
  NO2I1X1 g51827(.B (n_4482), .AN (n_6799), .Q (n_5012));
  NO2I1X1 g51828(.B (n_4459), .AN (n_6808), .Q (n_5011));
  NO2I1X1 g51829(.B (n_4490), .AN (n_6807), .Q (n_5010));
  NO2I1X1 g51830(.B (n_4753), .AN (n_6366), .Q (n_5009));
  NO2I1X1 g51831(.B (n_4753), .AN (n_6986), .Q (n_5008));
  NO2I1X1 g51832(.B (n_4459), .AN (n_6994), .Q (n_5007));
  NO2I1X1 g51833(.B (n_4747), .AN (n_6897), .Q (n_5006));
  NO2I1X1 g51834(.B (n_4485), .AN (n_6896), .Q (n_5005));
  NO2I1X1 g51835(.B (n_4742), .AN (n_6904), .Q (n_5004));
  NO2I1X1 g51836(.B (n_4743), .AN (n_6905), .Q (n_5003));
  NO2I1X1 g51837(.B (n_4747), .AN (n_6804), .Q (n_5002));
  NO2I1X1 g51838(.B (n_4486), .AN (n_6803), .Q (n_5001));
  NO2I1X1 g51839(.B (n_4743), .AN (n_6812), .Q (n_5000));
  NO2I1X1 g51840(.B (n_4742), .AN (n_6811), .Q (n_4999));
  AND2X1 g51841(.A (n_4741), .B (n_6784), .Q (n_4998));
  NO2I1X1 g51842(.B (n_4483), .AN (n_6350), .Q (n_4997));
  NO2I1X1 g51843(.B (n_4483), .AN (n_6970), .Q (n_4996));
  NO2I1X1 g51845(.B (n_4753), .AN (n_6304), .Q (n_4994));
  NO2I1X1 g51846(.B (n_4482), .AN (n_6303), .Q (n_4993));
  NO2I1X1 g51847(.B (n_4459), .AN (n_6312), .Q (n_4992));
  NO2I1X1 g51848(.B (n_4490), .AN (n_6311), .Q (n_4991));
  NO2I1X1 g51849(.B (n_4753), .AN (n_6273), .Q (n_4990));
  NO2I1X1 g51850(.B (n_4482), .AN (n_6272), .Q (n_4989));
  NO2I1X1 g51851(.B (n_4459), .AN (n_6281), .Q (n_4988));
  NO2I1X1 g51852(.B (n_4753), .AN (n_6552), .Q (n_4987));
  NO2I1X1 g51853(.B (n_4482), .AN (n_6551), .Q (n_4986));
  NO2I1X1 g51854(.B (n_4459), .AN (n_6560), .Q (n_4985));
  NO2I1X1 g51855(.B (n_4750), .AN (n_6559), .Q (n_4984));
  NO2I1X1 g51856(.B (n_4459), .AN (n_7118), .Q (n_4983));
  NO2I1X1 g51857(.B (n_4750), .AN (n_7117), .Q (n_4982));
  NO2I1X1 g51858(.B (n_4482), .AN (n_7109), .Q (n_4981));
  NO2I1X1 g51859(.B (n_4753), .AN (n_7110), .Q (n_4980));
  NO2I1X1 g51860(.B (n_4753), .AN (n_6397), .Q (n_4979));
  NO2I1X1 g51861(.B (n_4747), .AN (n_6308), .Q (n_4978));
  NO2I1X1 g51862(.B (n_4485), .AN (n_6307), .Q (n_4977));
  NO2I1X1 g51863(.B (n_4743), .AN (n_6316), .Q (n_4976));
  NO2I1X1 g51864(.B (n_4742), .AN (n_6315), .Q (n_4975));
  NO2I1X1 g51865(.B (n_4747), .AN (n_6277), .Q (n_4974));
  NO2I1X1 g51866(.B (n_4482), .AN (n_7202), .Q (n_4973));
  NO2I1X1 g51867(.B (n_4747), .AN (n_6556), .Q (n_4972));
  NO2I1X1 g51868(.B (n_4743), .AN (n_6564), .Q (n_4971));
  NO2I1X1 g51869(.B (n_4742), .AN (n_6563), .Q (n_4970));
  NO2I1X1 g51870(.B (n_4486), .AN (n_7113), .Q (n_4969));
  NO2I1X1 g51871(.B (n_4743), .AN (n_7122), .Q (n_4968));
  NO2I1X1 g51872(.B (n_4742), .AN (n_7121), .Q (n_4967));
  NO2I1X1 g51873(.B (n_4747), .AN (n_7114), .Q (n_4966));
  NO2I1X1 g51874(.B (n_4459), .AN (n_6932), .Q (n_4965));
  NO2I1X1 g51875(.B (n_4750), .AN (n_6931), .Q (n_4964));
  NO2I1X1 g51876(.B (n_4753), .AN (n_6924), .Q (n_4963));
  NO2I1X1 g51877(.B (n_4482), .AN (n_6923), .Q (n_4962));
  NO2I1X1 g51878(.B (n_4459), .AN (n_6870), .Q (n_4961));
  NO2I1X1 g51879(.B (n_4750), .AN (n_6869), .Q (n_4960));
  NO2I1X1 g51880(.B (n_4755), .AN (n_6862), .Q (n_4959));
  NO2I1X1 g51881(.B (n_4482), .AN (n_6861), .Q (n_4958));
  NO2I1X1 g51882(.B (n_4459), .AN (n_6839), .Q (n_4957));
  NO2I1X1 g51883(.B (n_4750), .AN (n_6838), .Q (n_4956));
  NO2I1X1 g51884(.B (n_4753), .AN (n_6831), .Q (n_4955));
  NO2I1X1 g51885(.B (n_4482), .AN (n_6830), .Q (n_4954));
  NO2I1X1 g51886(.B (n_4482), .AN (n_7078), .Q (n_4953));
  NO2I1X1 g51887(.B (n_4750), .AN (n_7179), .Q (n_4952));
  NO2I1X1 g51890(.B (n_4753), .AN (n_7141), .Q (n_4949));
  NO2I1X1 g51891(.B (n_4482), .AN (n_7140), .Q (n_4948));
  NO2I1X1 g51892(.B (n_4751), .AN (n_7148), .Q (n_4947));
  NO2I1X1 g51893(.B (n_4459), .AN (n_7149), .Q (n_4946));
  NO2I1X1 g51894(.B (n_4750), .AN (n_7086), .Q (n_4945));
  NO2I1X1 g51895(.B (n_4753), .AN (n_7079), .Q (n_4944));
  NO2I1X1 g51896(.B (n_4460), .AN (n_7017), .Q (n_4943));
  NO2I1X1 g51897(.B (n_4482), .AN (n_7016), .Q (n_4942));
  NO2I1X1 g51898(.B (n_4459), .AN (n_7025), .Q (n_4941));
  NO2I1X1 g51899(.B (n_4750), .AN (n_7024), .Q (n_4940));
  NO2I1X1 g51900(.B (n_4459), .AN (n_7087), .Q (n_4939));
  NO2I1X1 g51901(.B (n_4459), .AN (n_7180), .Q (n_4938));
  NO2I1X1 g51906(.B (n_4747), .AN (n_6928), .Q (n_4933));
  NO2I1X1 g51907(.B (n_4485), .AN (n_6927), .Q (n_4932));
  NO2I1X1 g51908(.B (n_4743), .AN (n_6936), .Q (n_4931));
  NO2I1X1 g51909(.B (n_4742), .AN (n_6935), .Q (n_4930));
  NO2I1X1 g51910(.B (n_4487), .AN (n_6866), .Q (n_4929));
  NO2I1X1 g51911(.B (n_4486), .AN (n_6865), .Q (n_4928));
  NO2I1X1 g51912(.B (n_4743), .AN (n_6874), .Q (n_4927));
  NO2I1X1 g51913(.B (n_4742), .AN (n_6873), .Q (n_4926));
  NO2I1X1 g51914(.B (n_4747), .AN (n_6835), .Q (n_4925));
  NO2I1X1 g51915(.B (n_4485), .AN (n_6834), .Q (n_4924));
  NO2I1X1 g51916(.B (n_4743), .AN (n_6843), .Q (n_4923));
  NO2I1X1 g51917(.B (n_4742), .AN (n_6842), .Q (n_4922));
  NO2I1X1 g51918(.B (n_4742), .AN (n_7090), .Q (n_4921));
  NO2I1X1 g51919(.B (n_4486), .AN (n_7175), .Q (n_4920));
  NO2I1X1 g51920(.B (n_4743), .AN (n_7184), .Q (n_4919));
  NO2I1X2 g51921(.B (n_4742), .AN (n_7183), .Q (n_4918));
  NO2I1X1 g51922(.B (n_4485), .AN (n_7144), .Q (n_4917));
  NO2I1X1 g51923(.B (n_4743), .AN (n_7153), .Q (n_4916));
  NO2I1X1 g51924(.B (n_4742), .AN (n_7152), .Q (n_4915));
  NO2I1X1 g51925(.B (n_4487), .AN (n_7145), .Q (n_4914));
  NO2I1X1 g51926(.B (n_4487), .AN (n_7176), .Q (n_4913));
  NO2I1X1 g51927(.B (n_4486), .AN (n_7082), .Q (n_4912));
  NO2I1X1 g51928(.B (n_4743), .AN (n_7091), .Q (n_4911));
  NO2I1X1 g51929(.B (n_4747), .AN (n_7083), .Q (n_4910));
  NO2I1X1 g51930(.B (n_4747), .AN (n_7021), .Q (n_4909));
  INX1 g51934(.A (n_4907), .Q (n_4906));
  INX1 g51935(.A (n_4905), .Q (n_4907));
  INX6 g51936(.A (n_4904), .Q (n_4903));
  INX8 g51937(.A (n_4902), .Q (n_4901));
  INX8 g51938(.A (n_4900), .Q (n_4899));
  INX6 g51939(.A (n_4898), .Q (n_4897));
  INX8 g51940(.A (n_4896), .Q (n_4895));
  INX6 g51941(.A (n_4894), .Q (n_4893));
  INX8 g51942(.A (n_4892), .Q (n_4891));
  BUX6 g51944(.A (n_4889), .Q (n_4888));
  INX1 g51946(.A (n_4888), .Q (n_4887));
  INX1 g51949(.A (n_4509), .Q (n_4886));
  INX8 g51951(.A (n_4885), .Q (n_4884));
  INX8 g51961(.A (n_4463), .Q (n_4508));
  INX2 g51968(.A (n_4883), .Q (n_4507));
  INX3 g51970(.A (n_4881), .Q (n_4882));
  INX2 g51972(.A (n_4883), .Q (n_4881));
  INX8 g51973(.A (n_4759), .Q (n_4883));
  INX8 g51979(.A (n_4880), .Q (n_4506));
  INX8 g51984(.A (n_4879), .Q (n_4878));
  INX4 g51989(.A (n_4877), .Q (n_4502));
  INX3 g51992(.A (n_4503), .Q (n_4877));
  BUX2 g51993(.A (n_4503), .Q (n_4876));
  INX4 g51998(.A (n_4452), .Q (n_4874));
  BUX3 g51999(.A (n_4452), .Q (n_4873));
  INX2 g52004(.A (n_4874), .Q (n_4500));
  INX8 g52007(.A (n_4871), .Q (n_4870));
  INX8 g52008(.A (n_4869), .Q (n_4868));
  INX6 g52010(.A (n_4865), .Q (n_4866));
  INX3 g52013(.A (n_4499), .Q (n_4865));
  BUX6 g52017(.A (n_4497), .Q (n_4498));
  INX6 g52019(.A (n_4457), .Q (n_4861));
  NO2I1X1 g52020(.B (n_4743), .AN (n_6688), .Q (n_4860));
  NO2I1X1 g52021(.B (n_4743), .AN (n_7029), .Q (n_4859));
  NO2I1X1 g52022(.B (n_4742), .AN (n_7028), .Q (n_4858));
  NO2I1X1 g52023(.B (n_4747), .AN (n_6339), .Q (n_4857));
  NO2I1X1 g52024(.B (n_4485), .AN (n_6338), .Q (n_4856));
  NO2I1X1 g52025(.B (n_4743), .AN (n_6347), .Q (n_4855));
  NO2I1X1 g52026(.B (n_4742), .AN (n_6346), .Q (n_4854));
  NO2I1X1 g52027(.B (n_4483), .AN (n_6257), .Q (n_4853));
  NO2I1X1 g52028(.B (n_4483), .AN (n_6536), .Q (n_4852));
  NO2I1X1 g52029(.B (n_4483), .AN (n_6381), .Q (n_4851));
  NO2I1X1 g52030(.B (n_4483), .AN (n_6288), .Q (n_4850));
  NO2I1X1 g52031(.B (n_4483), .AN (n_6846), .Q (n_4849));
  NO2I1X1 g52032(.B (n_4483), .AN (n_6815), .Q (n_4848));
  NO2I1X1 g52033(.B (n_4483), .AN (n_7156), .Q (n_4847));
  NO2I1X1 g52034(.B (n_4483), .AN (n_7125), .Q (n_4846));
  NO2I1X1 g52035(.B (n_4483), .AN (n_7063), .Q (n_4845));
  NO2I1X1 g52036(.B (n_4483), .AN (n_7001), .Q (n_4844));
  NO2I1X1 g52038(.B (n_4483), .AN (n_6908), .Q (n_4843));
  NO2I1X1 g52039(.B (n_4753), .AN (n_6769), .Q (n_4842));
  NO2I1X1 g52040(.B (n_4482), .AN (n_6768), .Q (n_4841));
  NO2I1X1 g52041(.B (n_4459), .AN (n_6777), .Q (n_4840));
  NO2I1X1 g52042(.B (n_4751), .AN (n_6776), .Q (n_4839));
  NO2I1X1 g52043(.B (n_4753), .AN (n_7048), .Q (n_4838));
  NO2I1X1 g52044(.B (n_4482), .AN (n_7047), .Q (n_4837));
  NO2I1X1 g52045(.B (n_4747), .AN (n_6773), .Q (n_4836));
  NO2I1X1 g52046(.B (n_4485), .AN (n_6772), .Q (n_4835));
  NO2I1X1 g52047(.B (n_4743), .AN (n_6781), .Q (n_4834));
  NO2I1X1 g52048(.B (n_4742), .AN (n_6780), .Q (n_4833));
  NO2I1X1 g52049(.B (n_4747), .AN (n_7052), .Q (n_4832));
  NO2I1X1 g52050(.B (n_4486), .AN (n_7051), .Q (n_4831));
  NO2I1X1 g52051(.B (n_4743), .AN (n_7060), .Q (n_4830));
  NO2I1X1 g52052(.B (n_4742), .AN (n_7059), .Q (n_4829));
  NA2X1 g52053(.A (n_4492), .B (n_6916), .Q (n_4828));
  NA2X1 g52054(.A (n_4478), .B (n_6915), .Q (n_4827));
  NO2I1X1 g52055(.B (n_4494), .AN (n_6823), .Q (n_4826));
  NO2I1X1 g52056(.B (n_4718), .AN (n_6822), .Q (n_4825));
  NO2I1X1 g52057(.B (n_4483), .AN (n_6753), .Q (n_4824));
  NO2I1X1 g52058(.B (n_4483), .AN (n_7032), .Q (n_4823));
  NA2X1 g52059(.A (n_4492), .B (n_7164), .Q (n_4822));
  NA2X1 g52060(.A (n_4478), .B (n_7163), .Q (n_4821));
  NO2I1X1 g52061(.B (n_4494), .AN (n_7071), .Q (n_4820));
  NO2I1X1 g52062(.B (n_4718), .AN (n_7070), .Q (n_4819));
  NO2I1X1 g52063(.B (n_4755), .AN (n_6738), .Q (n_4818));
  NO2I1X1 g52064(.B (n_4480), .AN (n_6737), .Q (n_4817));
  NO2I1X1 g52065(.B (n_4459), .AN (n_6746), .Q (n_4816));
  NO2I1X1 g52066(.B (n_4751), .AN (n_6745), .Q (n_4815));
  NO2I1X1 g52067(.B (n_4460), .AN (n_6707), .Q (n_4814));
  NO2I1X1 g52068(.B (n_4480), .AN (n_6706), .Q (n_4813));
  NO2I1X1 g52069(.B (n_4459), .AN (n_6715), .Q (n_4812));
  NO2I1X1 g52070(.B (n_4755), .AN (n_6676), .Q (n_4811));
  NO2I1X1 g52071(.B (n_4482), .AN (n_6675), .Q (n_4810));
  NO2I1X1 g52072(.B (n_4459), .AN (n_6684), .Q (n_4809));
  NO2I1X1 g52073(.B (n_4750), .AN (n_6683), .Q (n_4808));
  NO2I1X1 g52074(.B (n_4751), .AN (n_6714), .Q (n_4807));
  NO2I1X2 g52076(.B (n_4747), .AN (n_6742), .Q (n_4805));
  NO2I1X2 g52077(.B (n_4485), .AN (n_6741), .Q (n_4804));
  NO2I1X2 g52078(.B (n_4743), .AN (n_6750), .Q (n_4803));
  NO2I1X2 g52081(.B (n_4743), .AN (n_6719), .Q (n_4800));
  NO2I1X1 g52083(.B (n_4747), .AN (n_6680), .Q (n_4798));
  NO2I1X1 g52084(.B (n_4485), .AN (n_6679), .Q (n_4797));
  NO2I1X1 g52085(.B (n_4486), .AN (n_7020), .Q (n_4796));
  NO2I1X1 g52086(.B (n_4487), .AN (n_6711), .Q (n_4795));
  NO2I1X1 g52087(.B (n_4494), .AN (n_7040), .Q (n_4794));
  NO2I1X1 g52088(.B (n_4718), .AN (n_7039), .Q (n_4793));
  NA2X1 g52089(.A (n_4741), .B (n_6722), .Q (n_4792));
  NA2X1 g52090(.A (n_4741), .B (n_6691), .Q (n_4791));
  NA2X1 g52091(.A (n_4741), .B (n_6660), .Q (n_4790));
  NO2I1X1 g52093(.B (n_4718), .AN (n_6729), .Q (n_4789));
  NO2I1X1 g52094(.B (n_4483), .AN (n_6567), .Q (n_4788));
  NO2I1X1 g52095(.B (n_4459), .AN (n_6591), .Q (n_4787));
  NO2I1X1 g52096(.B (n_4486), .AN (n_6586), .Q (n_4786));
  NO2I1X1 g52097(.B (n_4487), .AN (n_6587), .Q (n_4785));
  NO2I1X1 g52098(.B (n_4460), .AN (n_6583), .Q (n_4784));
  NO2I1X1 g52099(.B (n_4480), .AN (n_6582), .Q (n_4783));
  NO2I1X2 g52100(.B (n_4490), .AN (n_6590), .Q (n_4782));
  NA2X1 g52101(.A (n_4741), .B (n_6629), .Q (n_4781));
  NO2I1X1 g52104(.B (n_4483), .AN (n_6474), .Q (n_4778));
  NA2X1 g52105(.A (n_4741), .B (n_6443), .Q (n_4777));
  AND2X1 g52106(.A (n_4488), .B (n_6463), .Q (n_4776));
  AND2X1 g52107(.A (n_4488), .B (n_6525), .Q (n_4775));
  AND2X1 g52108(.A (n_4488), .B (n_6618), .Q (n_4774));
  NO2I1X1 g52109(.B (n_4486), .AN (n_6617), .Q (n_4773));
  NO2I1X2 g52113(.B (n_4486), .AN (n_6524), .Q (n_4769));
  NO2I1X2 g52114(.B (n_4486), .AN (n_6462), .Q (n_4768));
  NA2X1 g52116(.A (n_4492), .B (n_6637), .Q (n_4766));
  NA2X1 g52117(.A (n_4478), .B (n_6636), .Q (n_4765));
  NA2X1 g52118(.A (n_4492), .B (n_6606), .Q (n_4764));
  NA2X1 g52119(.A (n_4478), .B (n_6605), .Q (n_4763));
  NA2X1 g52120(.A (n_4492), .B (n_6513), .Q (n_4762));
  NA2X1 g52121(.A (n_4478), .B (n_6512), .Q (n_4761));
  NO2I1X1 g52122(.B (n_4724), .AN (n_8480), .Q (n_8259));
  NO2I1X1 g52126(.B (n_4724), .AN (n_8484), .Q (n_8262));
  NA3X4 g52129(.A (n_4708), .B (n_4723), .C (n_4684), .Q (n_4908));
  NA2X2 g52130(.A (n_4723), .B (n_8482), .Q (n_4905));
  NA2X4 g52131(.A (n_4729), .B (n_4683), .Q (n_4904));
  NA2X4 g52132(.A (n_4729), .B (n_4694), .Q (n_4902));
  NA2X4 g52133(.A (n_4729), .B (n_4695), .Q (n_4900));
  NA2X4 g52134(.A (n_4730), .B (n_4695), .Q (n_4898));
  NA2X4 g52135(.A (n_4730), .B (n_4694), .Q (n_4896));
  NA2X4 g52136(.A (n_4730), .B (n_4683), .Q (n_4894));
  NA2X4 g52137(.A (n_4730), .B (n_4687), .Q (n_4892));
  NO2X4 g52138(.A (n_4688), .B (n_4726), .Q (n_4889));
  OR2X4 g52139(.A (n_4728), .B (n_4689), .Q (n_4885));
  NA2X4 g52141(.A (n_4727), .B (n_4695), .Q (n_4759));
  OR2X4 g52142(.A (n_4728), .B (n_4471), .Q (n_4880));
  OR2X4 g52143(.A (n_4726), .B (n_4682), .Q (n_4879));
  NA2I1X4 g52144(.B (n_4693), .AN (n_4728), .Q (n_4504));
  NO2I1X4 g52145(.B (n_4728), .AN (n_4693), .Q (n_4503));
  OR3X4 g52147(.A (n_4471), .B (n_4474), .C (n_4453), .Q (n_4871));
  OR3X4 g52148(.A (n_4471), .B (n_4477), .C (n_4453), .Q (n_4869));
  NO2X4 g52149(.A (n_4471), .B (n_4458), .Q (n_4499));
  OR2X4 g52150(.A (n_4471), .B (n_4458), .Q (n_4863));
  NO2X4 g52151(.A (n_4471), .B (n_4731), .Q (n_4497));
  OR2X4 g52152(.A (n_4471), .B (n_4731), .Q (n_4862));
  INX2 g52157(.A (n_4492), .Q (n_4494));
  BUX2 g52163(.A (n_4492), .Q (n_4756));
  BUX1 g52164(.A (n_4460), .Q (n_4755));
  INX6 g52165(.A (n_4752), .Q (n_4753));
  INX3 g52168(.A (n_4460), .Q (n_4752));
  INX2 g52171(.A (n_4489), .Q (n_4490));
  INX12 g52174(.A (n_4489), .Q (n_4751));
  BUX6 g52181(.A (n_4487), .Q (n_4747));
  BUX4 g52186(.A (n_4486), .Q (n_4485));
  INX6 g52189(.A (n_4744), .Q (n_4743));
  INX6 g52203(.A (n_4481), .Q (n_4482));
  INX3 g52204(.A (n_4740), .Q (n_4481));
  INX2 g52205(.A (n_4739), .Q (n_4740));
  INX1 g52207(.A (n_4739), .Q (n_4480));
  AND2X1 g52212(.A (n_4696), .B (instruction[28]), .Q (n_4737));
  AND2X1 g52213(.A (n_4696), .B (n_8480), .Q (n_4736));
  NA2X1 g52214(.A (n_4696), .B (n_8485), .Q (n_4735));
  NA2X1 g52215(.A (n_4696), .B (instruction[24]), .Q (n_4734));
  NA2X1 g52216(.A (n_4696), .B (n_8486), .Q (n_4733));
  AND2X1 g52217(.A (n_4696), .B (n_8481), .Q (n_4732));
  AND2X4 g52218(.A (n_4704), .B (n_4476), .Q (n_4492));
  NO2X2 g52220(.A (n_4707), .B (n_4474), .Q (n_4491));
  AND3X4 g52221(.A (n_4695), .B (n_4703), .C (n_4664), .Q (n_4489));
  NO2X2 g52222(.A (n_4707), .B (n_4701), .Q (n_4748));
  AND3X4 g52223(.A (n_4693), .B (n_4475), .C (n_4663), .Q (n_4488));
  NA2X4 g52224(.A (n_4706), .B (n_4475), .Q (n_4487));
  OR2X4 g52225(.A (n_4705), .B (n_4477), .Q (n_4486));
  NO2X4 g52226(.A (n_4705), .B (n_4477), .Q (n_4745));
  AND3X4 g52227(.A (n_4693), .B (n_4476), .C (n_4664), .Q (n_4744));
  AND3X4 g52228(.A (n_4693), .B (n_4703), .C (n_4663), .Q (n_4484));
  NA2X4 g52229(.A (n_4706), .B (n_4702), .Q (n_4742));
  AND2X4 g52230(.A (n_4704), .B (n_4475), .Q (n_4741));
  NA2X4 g52231(.A (n_4704), .B (n_4475), .Q (n_4483));
  NO2X4 g52232(.A (n_4707), .B (n_4477), .Q (n_4739));
  AND3X4 g52233(.A (n_4695), .B (n_4476), .C (n_4663), .Q (n_4738));
  INX1 g52235(.A (n_4728), .Q (n_4727));
  INX1 g52236(.A (n_4726), .Q (n_4725));
  INX4 g52237(.A (n_4724), .Q (n_4723));
  INX2 g52239(.A (n_4719), .Q (n_4720));
  INX2 g52240(.A (n_4478), .Q (n_4719));
  AND3X1 g52244(.A (n_4704), .B (n_4685), .C (n_4662), .Q (n_4717));
  AN22X1 g52245(.A (n_4692), .B (\instruction[10]_40063 ), .C (n_4472),
       .D (instruction[18]), .Q (n_4716));
  AN22X1 g52246(.A (n_4692), .B (\instruction[8]_40127 ), .C (n_4472),
       .D (n_4643), .Q (n_4715));
  AN22X1 g52247(.A (n_4692), .B (\instruction[9]_40095 ), .C (n_4472),
       .D (instruction[17]), .Q (n_4714));
  AN22X1 g52248(.A (n_4692), .B (\instruction[11]_40312 ), .C (n_4472),
       .D (n_4640), .Q (n_4713));
  AN22X1 g52249(.A (n_4472), .B (instruction[15]), .C (store_type), .D
       (\instruction[7]_39642 ), .Q (n_4712));
  NA2X1 g52250(.A (n_4696), .B (instruction[20]), .Q (n_4711));
  AN22X1 g52251(.A (branch_type), .B (\instruction[7]_39642 ), .C
       (jal_type), .D (instruction[20]), .Q (n_4710));
  NA2X4 g52252(.A (n_4698), .B (n_4664), .Q (n_4731));
  NO2X4 g52254(.A (n_4474), .B (n_4664), .Q (n_4730));
  NO2X4 g52255(.A (n_4477), .B (n_4664), .Q (n_4729));
  NA2X4 g52256(.A (n_4697), .B (n_4453), .Q (n_4728));
  NA2X4 g52257(.A (n_4699), .B (n_4453), .Q (n_4726));
  NA2I1X4 g52258(.B (n_4473), .AN (n_4696), .Q (n_4724));
  AND2X4 g52259(.A (n_4704), .B (n_4703), .Q (n_4478));
  NA2X2 g52260(.A (n_4704), .B (n_4702), .Q (n_4718));
  INX2 g52264(.A (n_4705), .Q (n_4706));
  AND2X2 g52266(.A (n_4691), .B (n_4473), .Q (n_4708));
  NA2X4 g52267(.A (n_4695), .B (n_4664), .Q (n_4707));
  NA2X4 g52268(.A (n_4693), .B (n_4663), .Q (n_4705));
  NO2X4 g52269(.A (n_4689), .B (n_4453), .Q (n_4704));
  INX1 g52272(.A (n_4701), .Q (n_4702));
  INX3 g52273(.A (n_4703), .Q (n_4701));
  INX2 g52274(.A (n_4700), .Q (n_4703));
  INX2 g52275(.A (n_4699), .Q (n_4700));
  BUX4 g52277(.A (n_4698), .Q (n_4476));
  BUX3 g52278(.A (n_4697), .Q (n_4698));
  INX3 g52280(.A (n_4474), .Q (n_4475));
  NA2X4 g52285(.A (n_4686), .B (n_4470), .Q (n_4477));
  NO2X2 g52286(.A (n_4686), .B (instruction[15]), .Q (n_4699));
  NO2I1X2 g52287(.B (n_4686), .AN (instruction[15]), .Q (n_4697));
  NA2X4 g52288(.A (n_4686), .B (instruction[15]), .Q (n_4474));
  NA2X4 g52289(.A (n_4690), .B (n_4680), .Q (n_4696));
  INX1 g52290(.A (n_4691), .Q (n_4692));
  BUX6 g52294(.A (n_4472), .Q (n_8157));
  INX1 g52295(.A (n_4473), .Q (n_4472));
  AND3X4 g52297(.A (n_4666), .B (n_8310), .C (n_4673), .Q (n_4695));
  NO2X4 g52298(.A (n_4677), .B (n_4666), .Q (n_4694));
  NO2I1X4 g52299(.B (n_4677), .AN (n_4675), .Q (n_4693));
  NO2X1 g52300(.A (branch_type), .B (n_4679), .Q (n_4691));
  INCX12 g52302(.A (n_4690), .Q (n_8296));
  INX3 g52305(.A (n_4689), .Q (n_4687));
  INX1 g52306(.A (n_4686), .Q (n_4685));
  INX1 g52307(.A (jal_type), .Q (n_4684));
  INX4 g52308(.A (n_4682), .Q (n_4683));
  NA2X2 g52311(.A (n_4678), .B (n_4668), .Q (n_4690));
  NA2X4 g52312(.A (n_4677), .B (n_4666), .Q (n_4689));
  NA2X4 g52313(.A (n_4667), .B (n_4676), .Q (n_4686));
  NO2X4 g52314(.A (n_8306), .B (n_8308), .Q (jal_type));
  NA2X4 g52315(.A (n_4677), .B (n_4675), .Q (n_4682));
  NA2X4 g52316(.A (n_4677), .B (n_4675), .Q (n_4471));
  INCX12 g52317(.A (n_4680), .Q (n_8166));
  BUX1 g52319(.A (n_4679), .Q (store_type));
  NA3I1X4 g52322(.B (n_4669), .C (n_4672), .AN (instruction[6]), .Q
       (n_4680));
  NO2I1X1 g52323(.B (n_4674), .AN (n_4670), .Q (system_type));
  NO3X2 g52324(.A (n_8302), .B (instruction[4]), .C (n_4661), .Q
       (n_4679));
  NO2X4 g52325(.A (n_4674), .B (n_8308), .Q (branch_type));
  INX1 g52326(.A (n_4678), .Q (n_8305));
  NA2X4 g52327(.A (n_4659), .B (n_4642), .Q (n_4676));
  NA2X1 g52328(.A (n_4672), .B (instruction[3]), .Q (n_8306));
  NO2X4 g52329(.A (n_4671), .B (instruction[3]), .Q (n_4678));
  INX4 g52331(.A (n_4666), .Q (n_4675));
  NA3X2 g52334(.A (instruction[1]), .B (n_4657), .C (instruction[0]),
       .Q (n_8302));
  NA3X4 g52335(.A (instruction[1]), .B (n_4656), .C (instruction[0]),
       .Q (n_4674));
  INX3 g52336(.A (n_4671), .Q (n_4672));
  NA2X4 g52337(.A (n_4667), .B (n_4640), .Q (n_4673));
  NA3X4 g52339(.A (instruction[1]), .B (instruction[0]), .C
       (instruction[2]), .Q (n_4671));
  INX1 g52340(.A (n_4669), .Q (n_8303));
  INX1 g52341(.A (n_4668), .Q (n_8304));
  NO2X1 g52342(.A (n_4658), .B (n_2416), .Q (n_8161));
  NO2X1 g52343(.A (n_4660), .B (n_4654), .Q (n_4670));
  NO2X4 g52344(.A (n_4661), .B (n_4654), .Q (n_4669));
  NO3X2 g52345(.A (n_4654), .B (instruction[6]), .C
       (\instruction[5]_40251 ), .Q (n_4668));
  BUX3 g52348(.A (n_4664), .Q (n_4663));
  MU2X1 g52350(.S (instruction[15]), .IN0 (n_6481), .IN1 (n_6482), .Q
       (n_4662));
  NO2X2 g52351(.A (n_4658), .B (\instruction[14]_40189 ), .Q (n_8163));
  NA3X2 g52352(.A (n_4644), .B (n_4641), .C (n_4639), .Q (n_4667));
  NA2X4 g52353(.A (n_4659), .B (n_4653), .Q (n_4666));
  NA2X4 g52355(.A (n_4655), .B (n_4646), .Q (n_4664));
  INX1 g52357(.A (n_4658), .Q (n_7302));
  NO2X1 g52358(.A (instruction[2]), .B (instruction[6]), .Q (n_4657));
  NO2X1 g52359(.A (instruction[2]), .B (n_4648), .Q (n_4656));
  NA2X2 g52360(.A (\instruction[5]_40251 ), .B (n_4649), .Q (n_4661));
  NA2X2 g52361(.A (instruction[6]), .B (\instruction[5]_40251 ), .Q
       (n_4660));
  NA2X4 g52362(.A (n_4644), .B (n_4639), .Q (n_4659));
  OR2X2 g52363(.A (n_8676), .B (n_8487), .Q (n_4658));
  INX4 g52365(.A (instruction[4]), .Q (n_4654));
  NA2X2 g52366(.A (n_4638), .B (n_4643), .Q (n_4655));
  NA2X4 g52367(.A (n_4645), .B (instruction[17]), .Q (n_4653));
  NO2X2 g52368(.A (n_4643), .B (n_4640), .Q (n_4652));
  AND2X1 g52369(.A (n_4641), .B (n_4639), .Q (n_4651));
  NA2X4 g52370(.A (n_4636), .B (n_4622), .Q (instruction[1]));
  NA2X4 g52371(.A (n_4637), .B (n_4631), .Q (instruction[0]));
  INX2 g52376(.A (n_4649), .Q (instruction[3]));
  AO22X1 g52378(.A (n_4468), .B (read_data[8]), .C (n_8224), .D
       (prev_instruction[8]), .Q (\instruction[8]_40127 ));
  AO22X1 g52379(.A (n_4468), .B (read_data[9]), .C (n_8224), .D
       (prev_instruction[9]), .Q (\instruction[9]_40095 ));
  AO22X1 g52380(.A (n_4468), .B (read_data[10]), .C (n_8224), .D
       (prev_instruction[10]), .Q (\instruction[10]_40063 ));
  AO22X1 g52381(.A (n_4468), .B (read_data[11]), .C (n_8224), .D
       (prev_instruction[11]), .Q (\instruction[11]_40312 ));
  AO22X1 g52383(.A (n_4468), .B (read_data[7]), .C (n_8224), .D
       (prev_instruction[7]), .Q (\instruction[7]_39642 ));
  NA2X2 g52384(.A (n_4620), .B (n_4613), .Q (instruction[28]));
  NA2X4 g52385(.A (n_4632), .B (n_4612), .Q (instruction[24]));
  NA2X4 g52389(.A (n_4630), .B (n_4614), .Q (\instruction[5]_40251 ));
  NA2X2 g52390(.A (n_4629), .B (n_4617), .Q (\instruction[14]_40189 ));
  NA2X4 g52391(.A (n_4633), .B (n_4615), .Q (instruction[2]));
  NA2X2 g52392(.A (n_4634), .B (n_4616), .Q (instruction[6]));
  NA2X2 g52393(.A (n_4628), .B (n_4611), .Q (n_4648));
  BUX4 g52396(.A (n_4645), .Q (n_4646));
  INX2 g52397(.A (n_4644), .Q (n_4645));
  BUX1 g52400(.A (n_4642), .Q (instruction[18]));
  INX2 g52401(.A (n_4641), .Q (n_4642));
  INX3 g52404(.A (n_4639), .Q (instruction[17]));
  INX2 g52410(.A (instruction[15]), .Q (n_4470));
  BUX4 g52411(.A (n_4638), .Q (instruction[15]));
  AN21X1 g52413(.A (n_4465), .B (prev_instruction[0]), .C
       (flush_37557), .Q (n_4637));
  AN21X1 g52414(.A (n_8224), .B (prev_instruction[1]), .C
       (flush_37557), .Q (n_4636));
  NA2X4 g52416(.A (n_4586), .B (n_4589), .Q (instruction[21]));
  NA2X4 g52417(.A (n_4599), .B (n_4595), .Q (instruction[23]));
  NA2X4 g52418(.A (n_4455), .B (n_4590), .Q (instruction[22]));
  NA2X4 g52422(.A (n_4587), .B (n_4588), .Q (instruction[20]));
  NO2X4 g52423(.A (n_4597), .B (n_4601), .Q (n_4644));
  NA2X4 g52424(.A (n_4593), .B (n_4598), .Q (n_4643));
  OA21X4 g52425(.A (n_4579), .B (n_6083), .C (n_4591), .Q (n_4641));
  NA2X4 g52426(.A (n_4594), .B (n_4454), .Q (n_4640));
  NO2X4 g52427(.A (n_4456), .B (n_4592), .Q (n_4639));
  NA2I1X4 g52428(.B (n_4596), .AN (n_4600), .Q (n_4638));
  NA2X2 g52430(.A (n_4467), .B (read_data[6]), .Q (n_4634));
  NA2X1 g52431(.A (n_4467), .B (read_data[2]), .Q (n_4633));
  NA2X1 g52432(.A (n_4467), .B (read_data[24]), .Q (n_4632));
  NA2X1 g52433(.A (n_4585), .B (read_data[0]), .Q (n_4631));
  NA2X1 g52434(.A (n_4585), .B (read_data[5]), .Q (n_4630));
  NA2X1 g52435(.A (n_4467), .B (read_data[14]), .Q (n_4629));
  NA2X1 g52436(.A (n_4585), .B (read_data[3]), .Q (n_4628));
  NA2X1 g52437(.A (n_4466), .B (read_data[4]), .Q (n_4627));
  NA2X1 g52442(.A (n_4467), .B (read_data[1]), .Q (n_4622));
  NA2X1 g52444(.A (n_4467), .B (read_data[28]), .Q (n_4620));
  NA2X1 g52447(.A (n_8224), .B (prev_instruction[14]), .Q (n_4617));
  NA2X1 g52448(.A (n_4465), .B (prev_instruction[6]), .Q (n_4616));
  NA2X1 g52449(.A (n_8224), .B (prev_instruction[2]), .Q (n_4615));
  NA2X1 g52450(.A (n_8224), .B (prev_instruction[5]), .Q (n_4614));
  NA2X1 g52451(.A (n_8224), .B (prev_instruction[28]), .Q (n_4613));
  NA2X1 g52452(.A (n_4465), .B (prev_instruction[24]), .Q (n_4612));
  NA2X1 g52453(.A (n_8224), .B (prev_instruction[3]), .Q (n_4611));
  NA2X1 g52456(.A (n_4465), .B (prev_instruction[4]), .Q (n_4608));
  NO2X2 g52463(.A (n_4579), .B (n_4572), .Q (n_4601));
  NO2I1X1 g52464(.B (n_4464), .AN (prev_instruction[15]), .Q (n_4600));
  NA2X2 g52466(.A (n_4465), .B (prev_instruction[23]), .Q (n_4599));
  NA2X1 g52467(.A (n_4581), .B (prev_instruction[16]), .Q (n_4598));
  NO2X2 g52468(.A (n_4584), .B (n_4567), .Q (n_4597));
  NA2X2 g52469(.A (n_4466), .B (read_data[15]), .Q (n_4596));
  NA2X1 g52470(.A (n_4469), .B (read_data[23]), .Q (n_4595));
  NA2X1 g52471(.A (n_4582), .B (read_data[19]), .Q (n_4594));
  NA2X1 g52472(.A (n_4469), .B (read_data[16]), .Q (n_4593));
  NO2I1X2 g52473(.B (n_4579), .AN (prev_instruction[17]), .Q (n_4592));
  NA2X1 g52475(.A (n_4582), .B (read_data[18]), .Q (n_4591));
  NA2X2 g52477(.A (n_4466), .B (read_data[22]), .Q (n_4590));
  NA2X2 g52478(.A (n_4469), .B (read_data[21]), .Q (n_4589));
  NA2X1 g52479(.A (n_4582), .B (read_data[20]), .Q (n_4588));
  NA2X2 g52480(.A (n_4581), .B (prev_instruction[20]), .Q (n_4587));
  NA2X2 g52481(.A (n_4581), .B (prev_instruction[21]), .Q (n_4586));
  BUX4 g52483(.A (n_4469), .Q (n_4585));
  BUX4 g52484(.A (n_4583), .Q (n_4469));
  BUX1 g52487(.A (n_4467), .Q (n_4468));
  BUX6 g52491(.A (n_4466), .Q (n_4467));
  INX4 g52492(.A (n_4584), .Q (n_4466));
  INX2 g52493(.A (n_4583), .Q (n_4584));
  NO2X4 g52495(.A (n_4578), .B (n_4575), .Q (n_4583));
  NO2X4 g52496(.A (n_4578), .B (n_4575), .Q (n_4582));
  INX8 g52498(.A (n_4580), .Q (n_8224));
  INX4 g52504(.A (n_4581), .Q (n_4580));
  BUX4 g52506(.A (n_4581), .Q (n_4465));
  INX6 g52507(.A (n_4464), .Q (n_4581));
  NA2X4 g52509(.A (n_4578), .B (n_4574), .Q (n_4464));
  NA2X4 g52510(.A (n_4578), .B (n_4576), .Q (n_4579));
  NA3X4 g52511(.A (n_4573), .B (n_4571), .C (n_4526), .Q (n_4578));
  ON21X2 g52512(.A (n_4526), .B (write_response), .C (n_4573), .Q
       (n_7714));
  INX4 g52516(.A (n_4575), .Q (n_4576));
  INX4 g52517(.A (n_4575), .Q (n_4574));
  NA2X4 g52518(.A (n_4568), .B (n_4570), .Q (n_4575));
  NO2X4 g52519(.A (n_4569), .B (halt), .Q (n_4573));
  NO2X1 g52520(.A (prev_instruction[16]), .B (prev_instruction[15]), .Q
       (n_4572));
  NA2X2 g52521(.A (prev_load_request), .B (read_response), .Q (n_4571));
  NO2X2 g52522(.A (current_state[3]), .B (current_state[2]), .Q
       (n_4570));
  NO2X4 g52523(.A (n_4527), .B (read_response), .Q (n_4569));
  NO2X4 g52525(.A (n_4528), .B (current_state[0]), .Q (n_4568));
  NO2X1 g52526(.A (read_data[16]), .B (read_data[15]), .Q (n_4567));
  INX1 g52527(.A (n_7188), .Q (n_4566));
  INX1 g52528(.A (n_7245), .Q (n_4565));
  INX1 g52529(.A (n_7192), .Q (n_4564));
  INX1 g52530(.A (n_7246), .Q (n_4563));
  INX1 g52531(.A (n_6521), .Q (n_4562));
  INX1 g52532(.A (n_6520), .Q (n_4561));
  INX1 g52533(.A (n_6615), .Q (n_4560));
  INX1 g52534(.A (n_6517), .Q (n_4559));
  INX1 g52535(.A (n_6614), .Q (n_4558));
  INX1 g52536(.A (n_6613), .Q (n_4557));
  INX1 g52537(.A (n_6516), .Q (n_4556));
  INX1 g52538(.A (n_6526), .Q (n_4555));
  INX1 g52539(.A (n_6619), .Q (n_4554));
  INX1 g52540(.A (n_6522), .Q (n_4553));
  INX1 g52541(.A (n_7050), .Q (n_4552));
  INX1 g52542(.A (n_6775), .Q (n_4551));
  INX1 g52543(.A (n_7054), .Q (n_4550));
  INX1 g52544(.A (n_6770), .Q (n_4549));
  INX1 g52545(.A (n_6758), .Q (n_4548));
  INX1 g52546(.A (n_6774), .Q (n_4547));
  INX1 g52547(.A (n_7055), .Q (n_4546));
  INX1 g52548(.A (n_6640), .Q (n_4545));
  INX1 g52549(.A (n_6760), .Q (n_4544));
  INX1 g52550(.A (n_6762), .Q (n_4543));
  INX1 g52551(.A (n_6763), .Q (n_4542));
  INX1 g52552(.A (n_6771), .Q (n_4541));
  INX1 g52553(.A (n_6756), .Q (n_4540));
  INX1 g52554(.A (n_6757), .Q (n_4539));
  INX1 g52555(.A (n_6754), .Q (n_4538));
  INX1 g52556(.A (n_7056), .Q (n_4537));
  INX1 g52557(.A (n_6761), .Q (n_4536));
  INX1 g52558(.A (n_6641), .Q (n_4535));
  INX1 g52559(.A (n_6650), .Q (n_4534));
  INX1 g52560(.A (n_6646), .Q (n_4533));
  INX1 g52561(.A (n_6459), .Q (n_4532));
  INX1 g52562(.A (n_6458), .Q (n_4531));
  INX1 g52563(.A (n_6460), .Q (n_4530));
  INX1 g52564(.A (n_6464), .Q (n_4529));
  INX2 g52565(.A (current_state[1]), .Q (n_4528));
  INX2 g52566(.A (n_8053), .Q (n_4527));
  INX4 g52569(.A (n_4576), .Q (flush_37557));
  NA2I1X4 g2(.B (n_4694), .AN (n_4726), .Q (n_4463));
  AND2X4 g52571(.A (n_4725), .B (n_4695), .Q (n_4452));
  NA2I1X2 g52572(.B (instruction[20]), .AN (n_4908), .Q (n_4462));
  NA2I1X4 g52574(.B (n_4475), .AN (n_4707), .Q (n_4460));
  NA2I1X4 g52575(.B (n_4476), .AN (n_4707), .Q (n_4459));
  NA2I1X4 g52576(.B (n_4664), .AN (n_4700), .Q (n_4458));
  NA2I1X4 g52577(.B (n_4729), .AN (n_4689), .Q (n_4457));
  NA3I1X4 g52578(.B (n_4670), .C (n_4658), .AN (n_4674), .Q (n_4473));
  NA2I1X4 g52579(.B (n_4654), .AN (n_4660), .Q (n_8308));
  AND2X4 g52580(.A (n_4655), .B (n_4646), .Q (n_4453));
  NA3I1X2 g52581(.B (n_4651), .C (n_4652), .AN (n_4638), .Q (n_8310));
  NA2I1X4 g52583(.B (prev_instruction[22]), .AN (n_4580), .Q (n_4455));
  NA2I1X2 g52584(.B (prev_instruction[19]), .AN (n_4579), .Q (n_4454));
  NA3I1X4 g52585(.B (n_4627), .C (n_4608), .AN (flush_37557), .Q
       (instruction[4]));
  INX2 g52595(.A (n_4889), .Q (n_4509));
  INX2 g52597(.A (n_4506), .Q (n_4505));
  NO2I1X1 g52599(.B (n_4904), .AN (n_6479), .Q (n_4510));
  AND2X1 g52601(.A (n_4473), .B (n_8482), .Q (n_8263));
  AND2X2 g52607(.A (n_5442), .B (n_5450), .Q (n_4517));
  AND2X1 g52611(.A (n_4723), .B (n_8481), .Q (n_8261));
  AND2X1 g52613(.A (n_4723), .B (instruction[28]), .Q (n_8260));
  AND2X1 g52629(.A (n_5634), .B (n_5615), .Q (n_4523));
  AND2X1 g52631(.A (n_5565), .B (n_5571), .Q (n_4522));
  NO2I1X1 g52633(.B (n_4457), .AN (n_6475), .Q (n_4511));
  AND6X1 g52635(.A (n_5924), .B (n_4523), .C (n_5719), .D (n_5727), .E
       (n_5698), .F (n_5706), .Q (n_4525));
  ON21X2 g52643(.A (n_5230), .B (n_2416), .C (n_5228), .Q (n_7688));
  AND2X2 g52645(.A (n_4582), .B (read_data[17]), .Q (n_4456));
  DFRQX1 \csr_mepc_reg[0] (.C (rc_gclk_199945), .D (n_4378), .Q
       (n_4431));
  DFRQX1 \csr_mepc_reg[1] (.C (rc_gclk_199945), .D (n_4380), .Q
       (n_4432));
  DFRQX1 csr_mip_meip_reg(.C (clock), .D (n_2551), .Q (n_4433));
  DFRX1 \csr_mip_mfip_reg[0] (.C (clock), .D (n_2557), .Q
       (UNCONNECTED), .QN (n_4436));
  DFRQX1 \csr_mip_mfip_reg[10] (.C (clock), .D (n_2550), .Q (n_4446));
  DFRQX1 \csr_mip_mfip_reg[11] (.C (clock), .D (n_2554), .Q (n_4447));
  DFRQX1 \csr_mip_mfip_reg[12] (.C (clock), .D (n_2549), .Q (n_4448));
  DFRQX1 \csr_mip_mfip_reg[13] (.C (clock), .D (n_2558), .Q (n_4449));
  DFRX1 \csr_mip_mfip_reg[14] (.C (clock), .D (n_2555), .Q
       (UNCONNECTED0), .QN (n_4450));
  DFRX1 \csr_mip_mfip_reg[15] (.C (clock), .D (n_2567), .Q
       (UNCONNECTED1), .QN (n_4451));
  DFRQX1 \csr_mip_mfip_reg[1] (.C (clock), .D (n_2562), .Q (n_4437));
  DFRQX1 \csr_mip_mfip_reg[2] (.C (clock), .D (n_2559), .Q (n_4438));
  DFRX1 \csr_mip_mfip_reg[3] (.C (clock), .D (n_2566), .Q
       (UNCONNECTED2), .QN (n_4439));
  DFRX1 \csr_mip_mfip_reg[4] (.C (clock), .D (n_2561), .Q
       (UNCONNECTED3), .QN (n_4440));
  DFRX1 \csr_mip_mfip_reg[5] (.C (clock), .D (n_2563), .Q
       (UNCONNECTED4), .QN (n_4441));
  DFRX1 \csr_mip_mfip_reg[6] (.C (clock), .D (n_2560), .Q
       (UNCONNECTED5), .QN (n_4442));
  DFRQX1 \csr_mip_mfip_reg[7] (.C (clock), .D (n_2564), .Q (n_4443));
  DFRX1 \csr_mip_mfip_reg[8] (.C (clock), .D (n_2553), .Q
       (UNCONNECTED6), .QN (n_4444));
  DFRQX1 \csr_mip_mfip_reg[9] (.C (clock), .D (n_2565), .Q (n_4445));
  DFRQX1 csr_mip_msip_reg(.C (clock), .D (n_2552), .Q (n_4435));
  DFRQX1 csr_mip_mtip_reg(.C (clock), .D (n_2556), .Q (n_4434));
  DFRQX1 \csr_utime_reg[0] (.C (clock), .D (real_time_clock[0]), .Q
       (csr_utime[0]));
  DFRQX1 \csr_utime_reg[10] (.C (clock), .D (real_time_clock[10]), .Q
       (csr_utime[10]));
  DFRX1 \csr_utime_reg[11] (.C (clock), .D (real_time_clock[11]), .Q
       (UNCONNECTED7), .QN (csr_utime[11]));
  DFRQX1 \csr_utime_reg[12] (.C (clock), .D (real_time_clock[12]), .Q
       (csr_utime[12]));
  DFRQX1 \csr_utime_reg[13] (.C (clock), .D (real_time_clock[13]), .Q
       (csr_utime[13]));
  DFRQX1 \csr_utime_reg[14] (.C (clock), .D (real_time_clock[14]), .Q
       (csr_utime[14]));
  DFRQX1 \csr_utime_reg[15] (.C (clock), .D (real_time_clock[15]), .Q
       (csr_utime[15]));
  DFRX1 \csr_utime_reg[16] (.C (clock), .D (real_time_clock[16]), .Q
       (UNCONNECTED8), .QN (csr_utime[16]));
  DFRQX1 \csr_utime_reg[17] (.C (clock), .D (real_time_clock[17]), .Q
       (csr_utime[17]));
  DFRQX1 \csr_utime_reg[18] (.C (clock), .D (real_time_clock[18]), .Q
       (csr_utime[18]));
  DFRX1 \csr_utime_reg[19] (.C (clock), .D (real_time_clock[19]), .Q
       (UNCONNECTED9), .QN (csr_utime[19]));
  DFRQX1 \csr_utime_reg[1] (.C (clock), .D (real_time_clock[1]), .Q
       (csr_utime[1]));
  DFRX1 \csr_utime_reg[20] (.C (clock), .D (real_time_clock[20]), .Q
       (UNCONNECTED10), .QN (csr_utime[20]));
  DFRX1 \csr_utime_reg[21] (.C (clock), .D (real_time_clock[21]), .Q
       (UNCONNECTED11), .QN (csr_utime[21]));
  DFRQX1 \csr_utime_reg[22] (.C (clock), .D (real_time_clock[22]), .Q
       (csr_utime[22]));
  DFRQX1 \csr_utime_reg[23] (.C (clock), .D (real_time_clock[23]), .Q
       (csr_utime[23]));
  DFRX1 \csr_utime_reg[24] (.C (clock), .D (real_time_clock[24]), .Q
       (UNCONNECTED12), .QN (csr_utime[24]));
  DFRQX1 \csr_utime_reg[25] (.C (clock), .D (real_time_clock[25]), .Q
       (csr_utime[25]));
  DFRQX1 \csr_utime_reg[26] (.C (clock), .D (real_time_clock[26]), .Q
       (csr_utime[26]));
  DFRQX1 \csr_utime_reg[27] (.C (clock), .D (real_time_clock[27]), .Q
       (csr_utime[27]));
  DFRQX1 \csr_utime_reg[28] (.C (clock), .D (real_time_clock[28]), .Q
       (csr_utime[28]));
  DFRQX1 \csr_utime_reg[29] (.C (clock), .D (real_time_clock[29]), .Q
       (csr_utime[29]));
  DFRQX1 \csr_utime_reg[2] (.C (clock), .D (real_time_clock[2]), .Q
       (csr_utime[2]));
  DFRQX1 \csr_utime_reg[30] (.C (clock), .D (real_time_clock[30]), .Q
       (csr_utime[30]));
  DFRX1 \csr_utime_reg[31] (.C (clock), .D (real_time_clock[31]), .Q
       (UNCONNECTED13), .QN (csr_utime[31]));
  DFRQX1 \csr_utime_reg[32] (.C (clock), .D (real_time_clock[32]), .Q
       (csr_utime[32]));
  DFRX1 \csr_utime_reg[33] (.C (clock), .D (real_time_clock[33]), .Q
       (UNCONNECTED14), .QN (csr_utime[33]));
  DFRX1 \csr_utime_reg[34] (.C (clock), .D (real_time_clock[34]), .Q
       (UNCONNECTED15), .QN (csr_utime[34]));
  DFRX1 \csr_utime_reg[35] (.C (clock), .D (real_time_clock[35]), .Q
       (UNCONNECTED16), .QN (csr_utime[35]));
  DFRQX1 \csr_utime_reg[36] (.C (clock), .D (real_time_clock[36]), .Q
       (csr_utime[36]));
  DFRQX1 \csr_utime_reg[37] (.C (clock), .D (real_time_clock[37]), .Q
       (csr_utime[37]));
  DFRQX1 \csr_utime_reg[38] (.C (clock), .D (real_time_clock[38]), .Q
       (csr_utime[38]));
  DFRX1 \csr_utime_reg[39] (.C (clock), .D (real_time_clock[39]), .Q
       (UNCONNECTED17), .QN (csr_utime[39]));
  DFRQX1 \csr_utime_reg[3] (.C (clock), .D (real_time_clock[3]), .Q
       (csr_utime[3]));
  DFRQX1 \csr_utime_reg[40] (.C (clock), .D (real_time_clock[40]), .Q
       (csr_utime[40]));
  DFRQX1 \csr_utime_reg[41] (.C (clock), .D (real_time_clock[41]), .Q
       (csr_utime[41]));
  DFRQX1 \csr_utime_reg[42] (.C (clock), .D (real_time_clock[42]), .Q
       (csr_utime[42]));
  DFRX1 \csr_utime_reg[43] (.C (clock), .D (real_time_clock[43]), .Q
       (UNCONNECTED18), .QN (csr_utime[43]));
  DFRQX1 \csr_utime_reg[44] (.C (clock), .D (real_time_clock[44]), .Q
       (csr_utime[44]));
  DFRQX1 \csr_utime_reg[45] (.C (clock), .D (real_time_clock[45]), .Q
       (csr_utime[45]));
  DFRQX1 \csr_utime_reg[46] (.C (clock), .D (real_time_clock[46]), .Q
       (csr_utime[46]));
  DFRQX1 \csr_utime_reg[47] (.C (clock), .D (real_time_clock[47]), .Q
       (csr_utime[47]));
  DFRX1 \csr_utime_reg[48] (.C (clock), .D (real_time_clock[48]), .Q
       (UNCONNECTED19), .QN (csr_utime[48]));
  DFRQX1 \csr_utime_reg[49] (.C (clock), .D (real_time_clock[49]), .Q
       (csr_utime[49]));
  DFRQX1 \csr_utime_reg[4] (.C (clock), .D (real_time_clock[4]), .Q
       (csr_utime[4]));
  DFRQX1 \csr_utime_reg[50] (.C (clock), .D (real_time_clock[50]), .Q
       (csr_utime[50]));
  DFRX1 \csr_utime_reg[51] (.C (clock), .D (real_time_clock[51]), .Q
       (UNCONNECTED20), .QN (csr_utime[51]));
  DFRX1 \csr_utime_reg[52] (.C (clock), .D (real_time_clock[52]), .Q
       (UNCONNECTED21), .QN (csr_utime[52]));
  DFRX1 \csr_utime_reg[53] (.C (clock), .D (real_time_clock[53]), .Q
       (UNCONNECTED22), .QN (csr_utime[53]));
  DFRQX1 \csr_utime_reg[54] (.C (clock), .D (real_time_clock[54]), .Q
       (csr_utime[54]));
  DFRQX1 \csr_utime_reg[55] (.C (clock), .D (real_time_clock[55]), .Q
       (csr_utime[55]));
  DFRX1 \csr_utime_reg[56] (.C (clock), .D (real_time_clock[56]), .Q
       (UNCONNECTED23), .QN (csr_utime[56]));
  DFRQX1 \csr_utime_reg[57] (.C (clock), .D (real_time_clock[57]), .Q
       (csr_utime[57]));
  DFRQX1 \csr_utime_reg[58] (.C (clock), .D (real_time_clock[58]), .Q
       (csr_utime[58]));
  DFRQX1 \csr_utime_reg[59] (.C (clock), .D (real_time_clock[59]), .Q
       (csr_utime[59]));
  DFRQX1 \csr_utime_reg[5] (.C (clock), .D (real_time_clock[5]), .Q
       (csr_utime[5]));
  DFRQX1 \csr_utime_reg[60] (.C (clock), .D (real_time_clock[60]), .Q
       (csr_utime[60]));
  DFRQX1 \csr_utime_reg[61] (.C (clock), .D (real_time_clock[61]), .Q
       (csr_utime[61]));
  DFRQX1 \csr_utime_reg[62] (.C (clock), .D (real_time_clock[62]), .Q
       (csr_utime[62]));
  DFRX1 \csr_utime_reg[63] (.C (clock), .D (real_time_clock[63]), .Q
       (UNCONNECTED24), .QN (csr_utime[63]));
  DFRQX1 \csr_utime_reg[6] (.C (clock), .D (real_time_clock[6]), .Q
       (csr_utime[6]));
  DFRX1 \csr_utime_reg[7] (.C (clock), .D (real_time_clock[7]), .Q
       (UNCONNECTED25), .QN (csr_utime[7]));
  DFRQX1 \csr_utime_reg[8] (.C (clock), .D (real_time_clock[8]), .Q
       (csr_utime[8]));
  DFRQX1 \csr_utime_reg[9] (.C (clock), .D (real_time_clock[9]), .Q
       (csr_utime[9]));
  DFRQX1 reset_reg_reg(.C (clock), .D (reset), .Q (reset_reg));
  AO22X2 g88822(.A (n_4381), .B (\instruction_address[0] ), .C
       (n_2309), .D (prev_rw_address[0]), .Q (n_7625));
  NA2X4 g88823(.A (n_4429), .B (n_8568), .Q (n_6235));
  NA2X4 g88824(.A (n_4430), .B (n_2718), .Q (n_7636));
  NA2X2 g88825(.A (n_4428), .B (n_4425), .Q (n_7304));
  NA2X2 g88826(.A (n_2719), .B (csr_data_out[0]), .Q (n_4430));
  ON31X1 g88827(.A (n_2507), .B (n_2585), .C (n_2583), .D
       (csr_data_out[1]), .Q (n_4429));
  ON21X1 g88828(.A (n_4424), .B (n_2297), .C (n_7882), .Q (n_4428));
  AO22X2 g88829(.A (n_4381), .B (n_8232), .C (n_2309), .D
       (prev_rw_address[1]), .Q (n_7626));
  AO22X1 g88831(.A (n_8231), .B (n_2475), .C
       (prev_instruction_address[0]), .D (n_2474), .Q
       (\instruction_address[0] ));
  NA3X1 g88832(.A (n_4426), .B (n_2975), .C (n_2971), .Q
       (csr_data_out[0]));
  NA3X2 g88833(.A (n_4427), .B (n_2926), .C (n_2924), .Q
       (csr_data_out[1]));
  AN221X1 g88834(.A (n_4432), .B (n_2323), .C (csr_mtval[1]), .D
       (n_2726), .E (n_8564), .Q (n_4427));
  AN221X1 g88835(.A (csr_mscratch[0]), .B (n_2727), .C (csr_mcause[0]),
       .D (n_2725), .E (n_4423), .Q (n_4426));
  AO22X1 g88836(.A (n_4396), .B (n_3203), .C (n_2309), .D
       (prev_write_strobe[2]), .Q (n_7631));
  AO22X1 g88837(.A (n_4396), .B (n_2278), .C (n_2309), .D
       (prev_write_strobe[3]), .Q (n_7628));
  NO3X2 g88838(.A (n_4422), .B (n_8216), .C (n_8222), .Q (n_4425));
  AO22X1 g88839(.A (n_4396), .B (n_3102), .C (n_2309), .D
       (prev_write_strobe[1]), .Q (n_7629));
  NA3X1 g88840(.A (n_4398), .B (n_4399), .C (n_4384), .Q (n_4424));
  AO22X1 g88841(.A (n_4396), .B (n_3110), .C (n_2309), .D
       (prev_write_strobe[0]), .Q (n_7630));
  AO222X2 g88842(.A (csr_utime[0]), .B (n_2619), .C (n_4431), .D
       (n_2729), .E (csr_utime[32]), .F (n_2312), .Q (n_4423));
  AO22X1 g88843(.A (n_960), .B (n_4431), .C (n_2386), .D
       (program_counter[0]), .Q (n_8231));
  ON21X1 g88844(.A (n_4363), .B (n_2628), .C (n_4421), .Q (n_8232));
  AO21X2 g88845(.A (n_4381), .B (n_8230), .C (n_4411), .Q (n_7619));
  AO21X2 g88846(.A (n_4381), .B (n_8233), .C (n_4415), .Q (n_7618));
  AO21X2 g88847(.A (n_4381), .B (n_8238), .C (n_4419), .Q (n_7613));
  AO21X2 g88848(.A (n_4381), .B (n_8237), .C (n_4418), .Q (n_7614));
  AO21X2 g88849(.A (n_4381), .B (n_8235), .C (n_4416), .Q (n_7616));
  AO21X2 g88850(.A (n_4381), .B (n_8236), .C (n_4417), .Q (n_7615));
  AO21X2 g88851(.A (n_4381), .B (n_8256), .C (n_4414), .Q (n_7627));
  AO21X2 g88852(.A (n_4381), .B (n_8234), .C (n_4412), .Q (n_7617));
  AO21X2 g88853(.A (n_4381), .B (n_8245), .C (n_4413), .Q (n_7606));
  AO21X2 g88854(.A (n_4381), .B (n_8225), .C (n_4406), .Q (n_7624));
  AO21X2 g88855(.A (n_4381), .B (n_8229), .C (n_4410), .Q (n_7620));
  AO21X2 g88856(.A (n_4381), .B (n_8228), .C (n_4409), .Q (n_7621));
  AO21X2 g88857(.A (n_4381), .B (n_8227), .C (n_4408), .Q (n_7622));
  AO21X2 g88858(.A (n_4381), .B (n_8226), .C (n_4407), .Q (n_7623));
  AO21X2 g88859(.A (n_4381), .B (n_8255), .C (n_4405), .Q (n_7596));
  AO21X2 g88860(.A (n_4381), .B (n_8254), .C (n_4404), .Q (n_7597));
  AO21X2 g88861(.A (n_4381), .B (n_8253), .C (n_4403), .Q (n_7598));
  AO21X2 g88862(.A (n_4381), .B (n_8252), .C (n_4402), .Q (n_7599));
  AO21X2 g88863(.A (n_4381), .B (n_8251), .C (n_4386), .Q (n_7600));
  AO21X2 g88864(.A (n_4381), .B (n_8240), .C (n_4387), .Q (n_7611));
  AO21X2 g88865(.A (n_4381), .B (n_8249), .C (n_4395), .Q (n_7602));
  AO21X2 g88866(.A (n_4381), .B (n_8248), .C (n_4394), .Q (n_7603));
  AO21X2 g88867(.A (n_4381), .B (n_8247), .C (n_4393), .Q (n_7604));
  AO21X2 g88868(.A (n_4381), .B (n_8246), .C (n_4392), .Q (n_7605));
  AO21X2 g88869(.A (n_4381), .B (n_8244), .C (n_4391), .Q (n_7607));
  AO21X2 g88870(.A (n_4381), .B (n_8243), .C (n_4390), .Q (n_7608));
  AO21X2 g88871(.A (n_4381), .B (n_8242), .C (n_4389), .Q (n_7609));
  AO21X2 g88872(.A (n_4381), .B (n_8241), .C (n_4388), .Q (n_7610));
  AO21X2 g88873(.A (n_4381), .B (n_8250), .C (n_4401), .Q (n_7601));
  AO21X2 g88874(.A (n_4381), .B (n_8239), .C (n_4420), .Q (n_7612));
  ON21X1 g88875(.A (n_4366), .B (n_2861), .C (n_4400), .Q (n_4422));
  NO2X1 g88876(.A (n_4397), .B (n_2810), .Q (n_8209));
  NO2X1 g88877(.A (n_4397), .B (n_2694), .Q (n_8211));
  NO2X1 g88878(.A (n_4397), .B (n_2693), .Q (n_8210));
  NO2X1 g88879(.A (n_4398), .B (n_2307), .Q (n_8214));
  NO2X1 g88880(.A (n_4399), .B (n_2307), .Q (n_8212));
  NA2X1 g88882(.A (n_960), .B (n_4432), .Q (n_4421));
  ON22X1 g88883(.A (n_2298), .B (n_2887), .C (n_8207), .D (n_6104), .Q
       (n_4420));
  ON22X1 g88884(.A (n_2298), .B (n_2916), .C (n_8207), .D (n_6105), .Q
       (n_4419));
  ON22X1 g88885(.A (n_2298), .B (n_2915), .C (n_8207), .D (n_6106), .Q
       (n_4418));
  ON22X1 g88886(.A (n_2298), .B (n_2914), .C (n_8207), .D (n_6107), .Q
       (n_4417));
  ON22X1 g88887(.A (n_2298), .B (n_2911), .C (n_8207), .D (n_6108), .Q
       (n_4416));
  ON22X1 g88888(.A (n_2298), .B (n_2912), .C (n_8207), .D (n_6111), .Q
       (n_4415));
  ON22X1 g88889(.A (n_2298), .B (n_2907), .C (n_8207), .D (n_6109), .Q
       (n_4414));
  ON22X1 g88890(.A (n_2298), .B (n_2906), .C (n_8207), .D (n_6110), .Q
       (n_4413));
  ON22X1 g88891(.A (n_2298), .B (n_2905), .C (n_8207), .D (n_6112), .Q
       (n_4412));
  ON22X1 g88892(.A (n_2298), .B (n_2904), .C (n_8207), .D (n_6113), .Q
       (n_4411));
  ON22X1 g88893(.A (n_2298), .B (n_2903), .C (n_8207), .D (n_6114), .Q
       (n_4410));
  ON22X1 g88894(.A (n_2298), .B (n_2902), .C (n_8207), .D (n_6085), .Q
       (n_4409));
  ON22X1 g88895(.A (n_2298), .B (n_2901), .C (n_8207), .D (n_6086), .Q
       (n_4408));
  ON22X1 g88896(.A (n_2298), .B (n_2910), .C (n_8207), .D (n_6087), .Q
       (n_4407));
  ON22X1 g88897(.A (n_2298), .B (n_2900), .C (n_8207), .D (n_6088), .Q
       (n_4406));
  ON22X1 g88898(.A (n_2298), .B (n_2899), .C (n_8207), .D (n_6089), .Q
       (n_4405));
  ON22X1 g88899(.A (n_2298), .B (n_2898), .C (n_8207), .D (n_6090), .Q
       (n_4404));
  ON22X1 g88900(.A (n_2298), .B (n_2908), .C (n_8207), .D (n_6091), .Q
       (n_4403));
  ON22X1 g88901(.A (n_2298), .B (n_2897), .C (n_8207), .D (n_6092), .Q
       (n_4402));
  ON22X1 g88902(.A (n_2298), .B (n_2909), .C (n_8207), .D (n_6094), .Q
       (n_4401));
  INX4 g88903(.A (n_2389), .Q (read_request));
  INX1 g88904(.A (n_8215), .Q (n_4400));
  BUCX4 g88905(.A (n_4396), .Q (write_request));
  ON22X1 g88906(.A (n_2298), .B (n_2896), .C (n_8207), .D (n_6095), .Q
       (n_4395));
  ON22X1 g88907(.A (n_2298), .B (n_2892), .C (n_8207), .D (n_6096), .Q
       (n_4394));
  ON22X1 g88908(.A (n_2298), .B (n_2890), .C (n_8207), .D (n_6097), .Q
       (n_4393));
  ON22X1 g88909(.A (n_2298), .B (n_2889), .C (n_8207), .D (n_6098), .Q
       (n_4392));
  ON22X1 g88910(.A (n_2298), .B (n_2891), .C (n_8207), .D (n_6099), .Q
       (n_4391));
  ON22X1 g88911(.A (n_2298), .B (n_2893), .C (n_8207), .D (n_6100), .Q
       (n_4390));
  ON22X1 g88912(.A (n_2298), .B (n_2895), .C (n_8207), .D (n_6101), .Q
       (n_4389));
  ON22X1 g88913(.A (n_2298), .B (n_2894), .C (n_8207), .D (n_6102), .Q
       (n_4388));
  ON22X1 g88914(.A (n_2298), .B (n_2888), .C (n_8207), .D (n_6103), .Q
       (n_4387));
  ON22X1 g88916(.A (n_2298), .B (n_2913), .C (n_8207), .D (n_6093), .Q
       (n_4386));
  NO2X1 g88917(.A (n_4384), .B (n_2307), .Q (n_8213));
  NO2X1 g88918(.A (n_4385), .B (n_2307), .Q (n_8217));
  NO2X4 g88919(.A (n_2388), .B (n_2814), .Q (n_8215));
  NA2X1 g88922(.A (n_4383), .B (n_2709), .Q (n_4399));
  NA2X1 g88923(.A (n_4382), .B (n_2809), .Q (n_4398));
  NO3X2 g88924(.A (n_2388), .B (n_2307), .C (n_2691), .Q (n_8216));
  NA2X1 g88925(.A (n_4383), .B (n_7882), .Q (n_4397));
  AO21X2 g88926(.A (n_4376), .B (n_2571), .C (n_2603), .Q (n_4396));
  INX4 g88950(.A (n_4377), .Q (n_4381));
  NO2X1 g88951(.A (n_4373), .B (n_2918), .Q (n_8220));
  AND3X1 g88959(.A (take_trap_39229), .B (program_counter[1]), .C
       (n_2503), .Q (n_4380));
  NA3X1 g88960(.A (n_4372), .B (n_2858), .C (n_2696), .Q (n_18082_BAR));
  NO2X1 g88961(.A (n_4373), .B (n_2807), .Q (n_8221));
  NO3X1 g88963(.A (n_4374), .B (n_4368), .C (n_4369), .Q (n_4379));
  NA2X1 g88964(.A (n_2279), .B (n_7882), .Q (n_18079_BAR));
  AND3X1 g88965(.A (take_trap_39229), .B (program_counter[0]), .C
       (n_2503), .Q (n_4378));
  NA2X1 g88966(.A (n_4375), .B (n_2503), .Q (n_7305));
  NA2X1 g88967(.A (n_4370), .B (n_2698), .Q (n_4385));
  NO3X2 g88968(.A (n_4373), .B (n_2759), .C (n_2692), .Q (n_8222));
  NA3X1 g88969(.A (n_4370), .B (n_2860), .C (n_2701), .Q (n_4384));
  NO2X1 g88970(.A (n_4371), .B (n_2947), .Q (n_4383));
  NO2X1 g88971(.A (n_4371), .B (n_2698), .Q (n_4382));
  AO21X2 g88972(.A (n_1169), .B (n_2945), .C (n_2570), .Q (n_4377));
  NA2X1 g88975(.A (n_1169), .B (n_2859), .Q (load_request_BAR));
  NA2X1 g88976(.A (n_4365), .B (n_7882), .Q (n_4375));
  AN31X1 g88977(.A (n_2697), .B (n_2695), .C (n_2763), .D (n_4367), .Q
       (n_4374));
  NO2X1 g88978(.A (take_trap_39229), .B (n_8569), .Q (n_4376));
  INX1 g88981(.A (n_4372), .Q (n_4373));
  INX1 g88982(.A (n_4371), .Q (n_4370));
  AND2X1 g88983(.A (n_4368), .B (n_7882), .Q (n_8223));
  NO2X1 g88984(.A (n_4366), .B (n_2762), .Q (n_8219));
  NO3X1 g88985(.A (n_4366), .B (n_2765), .C (n_2761), .Q (n_8218));
  NO2X1 g88987(.A (n_4367), .B (n_2307), .Q (n_4372));
  NA3I1X1 g88988(.B (n_4364), .C (n_7275), .AN (n_2984), .Q (n_4371));
  AO221X1 g88989(.A (n_7952), .B (n_2386), .C (n_4356), .D (n_7254), .E
       (n_2799), .Q (n_8229));
  AO221X1 g88990(.A (n_7929), .B (n_2386), .C (n_4356), .D (n_7273), .E
       (n_2751), .Q (n_8237));
  AO221X1 g88991(.A (n_7927), .B (n_2386), .C (n_4356), .D (n_7278), .E
       (n_2750), .Q (n_8236));
  AO221X1 g88992(.A (n_7926), .B (n_2386), .C (n_4356), .D (n_7279), .E
       (n_2749), .Q (n_8235));
  AO221X1 g88993(.A (n_7925), .B (n_2386), .C (n_4356), .D (n_7280), .E
       (n_2748), .Q (n_8233));
  AO221X1 g88994(.A (n_7956), .B (n_2386), .C (n_4356), .D (n_7251), .E
       (n_2796), .Q (n_8256));
  AO221X1 g88995(.A (n_7955), .B (n_2386), .C (n_4356), .D (n_7250), .E
       (n_2795), .Q (n_8245));
  AO221X1 g88996(.A (n_7954), .B (n_2386), .C (n_4356), .D (n_7252), .E
       (n_2794), .Q (n_8234));
  AO221X1 g88997(.A (n_7953), .B (n_2386), .C (n_4356), .D (n_7253), .E
       (n_2787), .Q (n_8230));
  AO221X1 g88998(.A (n_7930), .B (n_2386), .C (n_4356), .D (n_7272), .E
       (n_2752), .Q (n_8238));
  AO221X1 g88999(.A (n_7951), .B (n_2386), .C (n_4356), .D (n_7255), .E
       (n_2793), .Q (n_8228));
  AO221X1 g89000(.A (n_7950), .B (n_2386), .C (n_4356), .D (n_7256), .E
       (n_2792), .Q (n_8227));
  AO221X1 g89001(.A (n_7948), .B (n_2386), .C (n_4356), .D (n_7257), .E
       (n_2786), .Q (n_8226));
  AO221X1 g89002(.A (n_7947), .B (n_2386), .C (n_4356), .D (n_7258), .E
       (n_2798), .Q (n_8225));
  AO221X1 g89003(.A (n_7946), .B (n_2386), .C (n_4356), .D (n_7259), .E
       (n_2791), .Q (n_8255));
  AO221X1 g89004(.A (n_7945), .B (n_2386), .C (n_4356), .D (n_7260), .E
       (n_2790), .Q (n_8254));
  AO221X1 g89005(.A (n_7944), .B (n_2386), .C (n_4356), .D (n_7261), .E
       (n_2785), .Q (n_8253));
  AO221X1 g89006(.A (n_7943), .B (n_2386), .C (n_4356), .D (n_7262), .E
       (n_2797), .Q (n_8252));
  BUX12 g89012(.A (n_4365), .Q (take_trap_39229));
  NA2I1X1 g89013(.B (n_2780), .AN (n_4362), .Q (n_8184));
  NA2I1X1 g89014(.B (n_2779), .AN (n_4362), .Q (n_8204));
  NO2X1 g89015(.A (n_4361), .B (n_2760), .Q (n_4369));
  NO2X1 g89016(.A (n_4361), .B (n_2808), .Q (n_4368));
  AO221X1 g89017(.A (n_7938), .B (n_2386), .C (n_4356), .D (n_7268), .E
       (n_2801), .Q (n_8247));
  AO221X1 g89018(.A (n_7937), .B (n_2386), .C (n_4356), .D (n_7269), .E
       (n_2778), .Q (n_8246));
  AO221X1 g89019(.A (n_7936), .B (n_2386), .C (n_4356), .D (n_7277), .E
       (n_2772), .Q (n_8244));
  AO221X1 g89020(.A (n_7935), .B (n_2386), .C (n_4356), .D (n_7274), .E
       (n_2782), .Q (n_8243));
  AO221X1 g89021(.A (n_7934), .B (n_2386), .C (n_4356), .D (n_7270), .E
       (n_2777), .Q (n_8242));
  AO221X1 g89022(.A (n_7942), .B (n_2386), .C (n_4356), .D (n_7263), .E
       (n_2789), .Q (n_8251));
  AO221X1 g89023(.A (n_7932), .B (n_2386), .C (n_4356), .D (n_7266), .E
       (n_2754), .Q (n_8240));
  AO221X1 g89024(.A (n_7931), .B (n_2386), .C (n_4356), .D (n_7276), .E
       (n_2753), .Q (n_8239));
  AO221X1 g89025(.A (n_7933), .B (n_2386), .C (n_4356), .D (n_7271), .E
       (n_2771), .Q (n_8241));
  AO221X1 g89026(.A (n_7941), .B (n_2386), .C (n_4356), .D (n_7264), .E
       (n_2784), .Q (n_8250));
  NA2X1 g89027(.A (n_4364), .B (n_7275), .Q (n_4367));
  NA3X1 g89028(.A (n_4364), .B (n_2944), .C (n_7882), .Q (n_4366));
  AO221X1 g89029(.A (n_7940), .B (n_2386), .C (n_4356), .D (n_7265), .E
       (n_2781), .Q (n_8249));
  AO221X1 g89030(.A (n_7939), .B (n_2386), .C (n_4356), .D (n_7267), .E
       (n_2788), .Q (n_8248));
  NA2X4 g89031(.A (n_4360), .B (n_3384), .Q (n_4365));
  AN21X1 g89032(.A (n_2385), .B (program_counter[1]), .C (n_7862), .Q
       (n_4363));
  NO2X2 g89033(.A (n_4358), .B (n_4294), .Q (n_4364));
  INX1 g89034(.A (n_4360), .Q (n_4361));
  NA2X1 g89035(.A (n_4357), .B (n_4323), .Q (n_4362));
  NO2X2 g89036(.A (n_4358), .B (n_4241), .Q (n_4360));
  NO2X4 g89039(.A (n_4356), .B (n_2628), .Q (n_2386));
  BUX1 g89040(.A (n_4358), .Q (n_7862));
  NA2X1 g89041(.A (n_4356), .B (n_2964), .Q (n_4357));
  NO2X4 g89042(.A (n_2385), .B (n_957), .Q (n_4358));
  INX12 g89044(.A (n_2385), .Q (n_4356));
  NO2I1X4 g89049(.B (n_4355), .AN (n_2578), .Q (n_2385));
  NO2X2 g89050(.A (n_4354), .B (n_2500), .Q (n_4355));
  NO2X2 g89051(.A (n_4353), .B (n_4352), .Q (n_4354));
  ON21X1 g89052(.A (n_4350), .B (n_4313), .C (n_4349), .Q (n_4353));
  NA2X4 g89053(.A (n_4351), .B (n_4346), .Q (n_4352));
  NA2X2 g89054(.A (n_4350), .B (n_4314), .Q (n_4351));
  NO2X4 g89055(.A (n_4348), .B (n_4344), .Q (n_4350));
  NO2X2 g89056(.A (n_4347), .B (n_4285), .Q (n_4349));
  NO2X2 g89057(.A (n_4345), .B (n_2296), .Q (n_4348));
  NO2X4 g89058(.A (n_4343), .B (n_2418), .Q (n_4347));
  NA2X1 g89059(.A (n_4343), .B (n_8162), .Q (n_4346));
  NO2X2 g89060(.A (n_4342), .B (n_4339), .Q (n_4345));
  NA2X4 g89061(.A (n_4341), .B (n_4340), .Q (n_4344));
  NO2X2 g89062(.A (n_4338), .B (n_4328), .Q (n_4342));
  NA3X4 g89063(.A (n_4336), .B (n_4337), .C (n_4334), .Q (n_4343));
  NA2X2 g89064(.A (n_4335), .B (n_4316), .Q (n_4341));
  NO2X2 g89065(.A (n_4331), .B (n_4324), .Q (n_4340));
  NA2X2 g89066(.A (n_4332), .B (n_4330), .Q (n_4339));
  NO2X2 g89067(.A (n_4333), .B (n_4329), .Q (n_4338));
  NO2X2 g89068(.A (n_4328), .B (n_2293), .Q (n_4337));
  NO2X2 g89069(.A (n_4326), .B (n_4317), .Q (n_4336));
  NA2X2 g89070(.A (n_4325), .B (n_8489), .Q (n_4335));
  NO3X2 g89071(.A (n_2294), .B (n_4307), .C (n_4301), .Q (n_4334));
  NO2X2 g89072(.A (n_4319), .B (n_4277), .Q (n_4333));
  NA2X2 g89073(.A (n_4321), .B (n_4296), .Q (n_4332));
  NO2X2 g89074(.A (n_4320), .B (n_4295), .Q (n_4331));
  NO2X2 g89075(.A (n_4318), .B (n_2287), .Q (n_4330));
  NA2X2 g89076(.A (n_4322), .B (n_2290), .Q (n_4329));
  NA2X2 g89079(.A (n_4310), .B (n_4308), .Q (n_4326));
  NA2X2 g89080(.A (n_4312), .B (n_4306), .Q (n_4325));
  NA2X2 g89081(.A (n_4311), .B (n_4284), .Q (n_4324));
  NO2X1 g89082(.A (n_4315), .B (reset_internal_39074), .Q (n_4323));
  NA2X2 g89083(.A (n_4296), .B (n_4302), .Q (n_4328));
  NA2X1 g89084(.A (n_4297), .B (n_2383), .Q (n_4322));
  NA2X2 g89086(.A (n_4304), .B (n_2295), .Q (n_4321));
  NO2X2 g89087(.A (n_4303), .B (n_8653), .Q (n_4320));
  NO2X2 g89088(.A (n_4299), .B (n_4254), .Q (n_4319));
  NO2X2 g89089(.A (n_4298), .B (n_4252), .Q (n_4318));
  NA3X2 g89090(.A (n_4305), .B (n_4240), .C (n_4236), .Q (n_4317));
  AN21X1 g89092(.A (n_4242), .B (n_3384), .C (n_7714), .Q (n_4315));
  EO2X1 g89101(.A (alu_2nd_operand[11]), .B (alu_operation_code_39112),
       .Q (n_8284));
  AO21X1 g89102(.A (n_4240), .B (n_8161), .C (n_8159), .Q (n_4314));
  AN21X1 g89103(.A (n_4240), .B (n_8160), .C (n_8158), .Q (n_4313));
  EO2X1 g89105(.A (alu_2nd_operand[29]), .B (alu_operation_code_39112),
       .Q (n_8266));
  NA2X2 g89107(.A (n_4272), .B (n_4274), .Q (n_4312));
  NA2X2 g89108(.A (n_2286), .B (n_4250), .Q (n_4311));
  NO2X1 g89109(.A (n_4277), .B (n_4273), .Q (n_4310));
  MU2IX1 g89110(.S (alu_2nd_operand[28]), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8267));
  EO2X1 g89112(.A (alu_2nd_operand[27]), .B (alu_operation_code_39112),
       .Q (n_8268));
  NO3X1 g89116(.A (n_4262), .B (n_4230), .C (n_4245), .Q (n_4308));
  NA2X1 g89117(.A (n_2285), .B (n_2384), .Q (n_4307));
  NO2X1 g89118(.A (n_4278), .B (n_4177), .Q (n_4306));
  EO2X1 g89119(.A (alu_2nd_operand[31]), .B (alu_operation_code_39112),
       .Q (n_8264));
  NO2X2 g89122(.A (n_4295), .B (n_2292), .Q (n_4316));
  NO2X1 g89123(.A (n_2289), .B (n_4253), .Q (n_4305));
  MU2IX1 g89124(.S (alu_2nd_operand[15]), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8280));
  NA2X1 g89125(.A (n_4267), .B (n_4255), .Q (n_8289));
  MU2X1 g89126(.S (alu_2nd_operand[7]), .IN0
       (alu_operation_code_39112), .IN1 (n_2326), .Q (n_8288));
  EN2X1 g89127(.A (alu_2nd_operand[10]), .B (n_2326), .Q (n_8285));
  NA2X2 g89128(.A (n_4268), .B (n_2376), .Q (n_4304));
  EN2X1 g89129(.A (alu_2nd_operand[9]), .B (n_2326), .Q (n_8286));
  MU2IX1 g89130(.S (alu_2nd_operand[8]), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8287));
  NO2X1 g89131(.A (n_4256), .B (n_4244), .Q (n_4303));
  NO2X1 g89133(.A (n_4279), .B (n_4162), .Q (n_4302));
  MU2X1 g89134(.S (alu_2nd_operand[24]), .IN0
       (alu_operation_code_39112), .IN1 (n_2326), .Q (n_8271));
  MU2X1 g89135(.S (alu_2nd_operand[19]), .IN0
       (alu_operation_code_39112), .IN1 (n_2326), .Q (n_8276));
  NA3I1X2 g89136(.B (n_4213), .C (n_4228), .AN (n_2284), .Q (n_4301));
  MU2IX1 g89137(.S (alu_2nd_operand[25]), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8270));
  EN2X1 g89139(.A (n_8317), .B (n_2326), .Q (n_8265));
  EN2X1 g89140(.A (alu_2nd_operand[22]), .B (n_2326), .Q (n_8273));
  EN2X1 g89141(.A (alu_2nd_operand[21]), .B (n_2326), .Q (n_8274));
  MU2IX1 g89142(.S (alu_2nd_operand[26]), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8269));
  MU2IX1 g89144(.S (alu_2nd_operand[23]), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8272));
  MU2X1 g89145(.S (alu_2nd_operand[12]), .IN0
       (alu_operation_code_39112), .IN1 (n_2326), .Q (n_8283));
  NO3X2 g89147(.A (n_4227), .B (n_4214), .C (n_2374), .Q (n_4299));
  NO2X1 g89148(.A (n_4263), .B (n_2382), .Q (n_4298));
  NA2X1 g89149(.A (n_4270), .B (n_4212), .Q (n_4297));
  MU2IX1 g89151(.S (alu_2nd_operand[3]), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8292));
  MU2IX1 g89152(.S (n_8499), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8295));
  MU2IX1 g89153(.S (alu_2nd_operand[1]), .IN0 (n_2326), .IN1
       (alu_operation_code_39112), .Q (n_8294));
  NA3X1 g89154(.A (n_4242), .B (n_2760), .C (n_2700), .Q (n_4294));
  AO222X2 g89155(.A (n_2316), .B (n_4129), .C (n_2364), .D (n_3109), .E
       (prev_write_data[23]), .F (n_2309), .Q (write_data[23]));
  AO222X2 g89156(.A (n_2316), .B (n_2368), .C (n_2362), .D (n_3109), .E
       (prev_write_data[22]), .F (n_2309), .Q (write_data[22]));
  AO222X2 g89157(.A (n_2316), .B (n_2371), .C (n_2367), .D (n_3109), .E
       (prev_write_data[20]), .F (n_2309), .Q (write_data[20]));
  AO222X2 g89158(.A (n_2316), .B (n_4142), .C (n_4118), .D (n_3109), .E
       (prev_write_data[19]), .F (n_2309), .Q (write_data[19]));
  AO222X2 g89159(.A (n_2316), .B (n_4154), .C (n_4124), .D (n_3109), .E
       (prev_write_data[18]), .F (n_2309), .Q (write_data[18]));
  AO222X2 g89160(.A (n_2316), .B (n_4144), .C (n_4119), .D (n_3109), .E
       (prev_write_data[17]), .F (n_2309), .Q (write_data[17]));
  AO222X2 g89161(.A (n_2316), .B (n_4147), .C (n_8501), .D (n_3109), .E
       (prev_write_data[16]), .F (n_2309), .Q (write_data[16]));
  AO222X2 g89162(.A (n_2316), .B (n_2370), .C (n_4130), .D (n_3109), .E
       (prev_write_data[21]), .F (n_2309), .Q (write_data[21]));
  AO222X2 g89163(.A (n_4133), .B (n_3042), .C (n_2364), .D (n_3043), .E
       (prev_write_data[15]), .F (n_2309), .Q (write_data[15]));
  AO222X2 g89164(.A (n_4138), .B (n_3042), .C (n_2362), .D (n_3043), .E
       (prev_write_data[14]), .F (n_2309), .Q (write_data[14]));
  AO222X2 g89165(.A (n_4132), .B (n_3042), .C (n_4130), .D (n_3043), .E
       (prev_write_data[13]), .F (n_2309), .Q (write_data[13]));
  AO222X2 g89166(.A (n_4125), .B (n_3042), .C (n_4124), .D (n_3043), .E
       (prev_write_data[10]), .F (n_2309), .Q (write_data[10]));
  AO222X2 g89167(.A (n_4128), .B (n_3042), .C (n_4118), .D (n_3043), .E
       (prev_write_data[11]), .F (n_2309), .Q (write_data[11]));
  AO222X2 g89168(.A (n_4135), .B (n_3042), .C (n_8501), .D (n_3043), .E
       (prev_write_data[8]), .F (n_2309), .Q (write_data[8]));
  AO222X2 g89169(.A (n_4126), .B (n_3042), .C (n_2367), .D (n_3043), .E
       (prev_write_data[12]), .F (n_2309), .Q (write_data[12]));
  AO222X2 g89170(.A (n_4127), .B (n_3042), .C (n_4119), .D (n_3043), .E
       (prev_write_data[9]), .F (n_2309), .Q (write_data[9]));
  AN222X0 g89171(.A (n_2316), .B (n_4149), .C (prev_write_data[31]), .D
       (n_2309), .E (n_2968), .F (n_4133), .Q (n_4293));
  AN222X1 g89172(.A (n_2316), .B (n_4151), .C (prev_write_data[30]), .D
       (n_2309), .E (n_2968), .F (n_4138), .Q (n_4292));
  AN222X1 g89173(.A (n_2316), .B (n_4152), .C (prev_write_data[29]), .D
       (n_2309), .E (n_2968), .F (n_4132), .Q (n_4291));
  AN222X0 g89174(.A (n_2316), .B (n_4150), .C (prev_write_data[28]), .D
       (n_2309), .E (n_2968), .F (n_4126), .Q (n_4290));
  AN222X0 g89175(.A (n_2316), .B (n_4137), .C (prev_write_data[27]), .D
       (n_2309), .E (n_2968), .F (n_4128), .Q (n_4289));
  AN222X0 g89176(.A (n_2316), .B (n_8619), .C (prev_write_data[26]), .D
       (n_2309), .E (n_2968), .F (n_4125), .Q (n_4288));
  AN222X0 g89177(.A (n_2316), .B (n_4145), .C (prev_write_data[25]), .D
       (n_2309), .E (n_2968), .F (n_4127), .Q (n_4287));
  AN222X0 g89178(.A (n_2316), .B (n_4140), .C (prev_write_data[24]), .D
       (n_2309), .E (n_2968), .F (n_4135), .Q (n_4286));
  NO2X1 g89179(.A (n_4240), .B (n_2680), .Q (n_4285));
  ON21X1 g89180(.A (n_4203), .B (n_4208), .C (n_4200), .Q (n_4284));
  NO2X2 g89186(.A (n_4231), .B (n_4252), .Q (n_4296));
  NA2X2 g89187(.A (n_4250), .B (n_2384), .Q (n_4295));
  NA2X1 g89195(.A (n_4249), .B (n_4174), .Q (n_4274));
  NA2X1 g89196(.A (n_4251), .B (n_4246), .Q (n_4273));
  NO2X1 g89197(.A (n_4237), .B (n_8493), .Q (n_4272));
  ON21X1 g89199(.A (n_2373), .B (n_2306), .C (n_4131), .Q (n_4270));
  NA2X2 g89202(.A (n_4228), .B (n_4234), .Q (n_4268));
  NA2X1 g89203(.A (alu_2nd_operand[6]), .B (n_2326), .Q (n_4267));
  AN21X1 g89206(.A (n_2380), .B (n_4172), .C (n_2381), .Q (n_4264));
  NO2X1 g89207(.A (n_4215), .B (n_4132), .Q (n_4263));
  NA3X1 g89208(.A (n_4210), .B (n_2283), .C (n_2372), .Q (n_4262));
  AN21X1 g89217(.A (n_4178), .B (n_4179), .C (n_4176), .Q (n_4256));
  NA2X1 g89218(.A (n_4221), .B (alu_operation_code_39112), .Q (n_4255));
  NA2X1 g89219(.A (n_4239), .B (n_4175), .Q (n_4254));
  NA3I1X1 g89220(.B (n_2267), .C (n_4173), .AN (n_2374), .Q (n_4253));
  NA3X2 g89221(.A (n_2376), .B (n_4182), .C (n_2273), .Q (n_4279));
  NA2I1X4 g89222(.B (n_4235), .AN (n_4247), .Q (n_4278));
  NA2X1 g89223(.A (n_2383), .B (n_8494), .Q (n_4277));
  INX1 g89228(.A (n_4243), .Q (alu_2nd_operand[14]));
  INX1 g89229(.A (n_4241), .Q (n_4242));
  NA2X1 g89230(.A (n_2378), .B (n_2272), .Q (n_4239));
  AO22X4 g89231(.A (n_3110), .B (n_2367), .C (n_2309), .D
       (prev_write_data[4]), .Q (write_data[4]));
  AO22X4 g89232(.A (n_3110), .B (n_4118), .C (n_2309), .D
       (prev_write_data[3]), .Q (write_data[3]));
  AO22X4 g89233(.A (n_3110), .B (n_4124), .C (n_2309), .D
       (prev_write_data[2]), .Q (write_data[2]));
  AO22X4 g89234(.A (n_3110), .B (n_8501), .C (n_2309), .D
       (prev_write_data[0]), .Q (write_data[0]));
  AO22X4 g89235(.A (n_3110), .B (n_4130), .C (n_2309), .D
       (prev_write_data[5]), .Q (write_data[5]));
  AO22X4 g89236(.A (n_3110), .B (n_4119), .C (n_2309), .D
       (prev_write_data[1]), .Q (write_data[1]));
  AO22X4 g89237(.A (n_3110), .B (n_2364), .C (n_2309), .D
       (prev_write_data[7]), .Q (write_data[7]));
  NA2X1 g89238(.A (n_4202), .B (n_2269), .Q (n_4238));
  AO22X4 g89239(.A (n_3110), .B (n_2362), .C (n_2309), .D
       (prev_write_data[6]), .Q (write_data[6]));
  NO2X1 g89240(.A (n_4207), .B (n_4206), .Q (n_4237));
  NO2X1 g89241(.A (n_4202), .B (n_4189), .Q (n_4236));
  NO2X1 g89242(.A (n_4186), .B (n_4171), .Q (n_4235));
  NA2X1 g89243(.A (n_2377), .B (n_4182), .Q (n_4234));
  NO2X1 g89245(.A (n_4177), .B (n_4166), .Q (n_4232));
  NA2X1 g89246(.A (n_2265), .B (n_4159), .Q (n_4231));
  OR2X2 g89247(.A (n_4176), .B (n_4178), .Q (n_4230));
  NA2X1 g89248(.A (n_2379), .B (n_6135), .Q (n_4229));
  NA2X2 g89250(.A (n_4193), .B (n_4205), .Q (n_4252));
  NO2X2 g89252(.A (n_4195), .B (n_4190), .Q (n_4251));
  AND2X4 g89253(.A (n_4200), .B (n_2267), .Q (n_4250));
  NO2X2 g89254(.A (n_4206), .B (n_4185), .Q (n_4249));
  NA2X2 g89256(.A (n_4180), .B (n_2274), .Q (n_4247));
  NO2X1 g89257(.A (n_4194), .B (n_4156), .Q (n_4246));
  NA2X2 g89258(.A (n_4179), .B (n_4165), .Q (n_4245));
  NA2X2 g89259(.A (n_4198), .B (n_2472), .Q (alu_2nd_operand[13]));
  NA2X1 g89260(.A (n_4187), .B (n_4161), .Q (n_4244));
  MU2X2 g89261(.S (n_2258), .IN0 (n_7672), .IN1 (n_4152), .Q
       (alu_2nd_operand[29]));
  MU2IX1 g89262(.S (n_2258), .IN0 (n_7688), .IN1 (n_4138), .Q (n_4243));
  MU2X1 g89263(.S (n_2258), .IN0 (n_7673), .IN1 (n_4150), .Q
       (alu_2nd_operand[28]));
  MU2X1 g89264(.S (n_2258), .IN0 (n_8263), .IN1 (n_4149), .Q
       (alu_2nd_operand[31]));
  OR2X2 g89265(.A (n_8297), .B (n_4169), .Q (n_4241));
  NO2X2 g89266(.A (n_4199), .B (n_4203), .Q (n_4240));
  INX1 g89268(.A (n_4225), .Q (alu_2nd_operand[5]));
  INX1 g89269(.A (n_4224), .Q (alu_2nd_operand[17]));
  INX2 g89270(.A (n_4223), .Q (alu_2nd_operand[20]));
  INX1 g89272(.A (n_4221), .Q (alu_2nd_operand[6]));
  INX3 g89274(.A (n_8496), .Q (alu_2nd_operand[2]));
  INX1 g89275(.A (n_8497), .Q (alu_2nd_operand[18]));
  INX4 g89278(.A (n_828), .Q (alu_2nd_operand[1]));
  BUX8 g89279(.A (n_8499), .Q (alu_2nd_operand[0]));
  NO2X1 g89281(.A (n_4170), .B (\rs1_data[13]_39536 ), .Q (n_4215));
  NO2X1 g89282(.A (n_4173), .B (n_2375), .Q (n_4214));
  AN21X1 g89283(.A (n_4116), .B (n_6121), .C (n_2377), .Q (n_4213));
  NA2X1 g89284(.A (n_2373), .B (n_2306), .Q (n_4212));
  AN21X1 g89287(.A (n_4131), .B (n_2306), .C (n_2373), .Q (n_4210));
  NO2X2 g89288(.A (n_4197), .B (n_4155), .Q (n_4228));
  NA2X1 g89289(.A (n_2271), .B (n_4167), .Q (n_4227));
  NO2X1 g89290(.A (n_4196), .B (n_4164), .Q (n_4226));
  OA22X1 g89291(.A (n_4131), .B (n_2303), .C (n_2457), .D (n_2258), .Q
       (n_4225));
  OA22X1 g89292(.A (n_4143), .B (n_2303), .C (n_2462), .D (n_2258), .Q
       (n_4224));
  OA22X2 g89293(.A (n_4148), .B (n_2303), .C (n_2459), .D (n_2258), .Q
       (n_4223));
  MU2IX2 g89294(.S (n_2258), .IN0 (n_2458), .IN1 (n_4134), .Q
       (alu_2nd_operand[8]));
  MU2IX2 g89296(.S (n_2258), .IN0 (n_2460), .IN1 (n_2369), .Q
       (alu_2nd_operand[21]));
  MU2X2 g89297(.S (n_2258), .IN0 (n_7675), .IN1 (n_8619), .Q
       (alu_2nd_operand[26]));
  MU2X2 g89298(.S (n_2258), .IN0 (n_7691), .IN1 (n_4128), .Q
       (alu_2nd_operand[11]));
  MU2X2 g89299(.S (n_2258), .IN0 (n_7676), .IN1 (n_4145), .Q
       (alu_2nd_operand[25]));
  MU2X2 g89301(.S (n_2258), .IN0 (n_7683), .IN1 (n_4142), .Q
       (alu_2nd_operand[19]));
  MU2X1 g89302(.S (n_2258), .IN0 (n_8259), .IN1 (n_2363), .Q
       (alu_2nd_operand[7]));
  MU2IX1 g89303(.S (n_2258), .IN0 (n_8258), .IN1 (n_2362), .Q (n_4221));
  MU2X4 g89304(.S (n_2258), .IN0 (n_7677), .IN1 (n_4140), .Q
       (alu_2nd_operand[24]));
  MU2X1 g89305(.S (n_2258), .IN0 (n_7678), .IN1 (n_4129), .Q
       (alu_2nd_operand[23]));
  MU2X2 g89306(.S (n_2258), .IN0 (n_7687), .IN1 (n_4133), .Q
       (alu_2nd_operand[15]));
  MU2X2 g89307(.S (n_2258), .IN0 (n_8261), .IN1 (n_4127), .Q
       (alu_2nd_operand[9]));
  MU2X1 g89310(.S (n_2258), .IN0 (n_8262), .IN1 (n_4125), .Q
       (alu_2nd_operand[10]));
  MU2X4 g89311(.S (n_2258), .IN0 (n_7674), .IN1 (n_4137), .Q
       (alu_2nd_operand[27]));
  MU2X4 g89312(.S (n_2258), .IN0 (n_7690), .IN1 (n_4126), .Q
       (alu_2nd_operand[12]));
  MU2X4 g89313(.S (n_2258), .IN0 (n_7680), .IN1 (n_4118), .Q
       (alu_2nd_operand[3]));
  OA22X4 g89315(.A (n_2366), .B (n_2303), .C (n_2439), .D (n_2258), .Q
       (n_828));
  INX1 g89325(.A (n_4200), .Q (n_4199));
  NA2X2 g89327(.A (n_4132), .B (n_2258), .Q (n_4198));
  NO2I1X1 g89329(.B (n_4128), .AN (\rs1_data[11]_39506 ), .Q (n_4197));
  NO2I1X1 g89330(.B (n_2363), .AN (\rs1_data[7]_39466 ), .Q (n_4196));
  NO2I1X1 g89332(.B (n_4138), .AN (\rs1_data[14]_39546 ), .Q (n_4195));
  NO2I1X1 g89333(.B (n_2368), .AN (\rs1_data[22]_39626 ), .Q (n_4194));
  NA2X1 g89334(.A (n_4138), .B (n_2425), .Q (n_4193));
  NA2X1 g89335(.A (n_2362), .B (n_2428), .Q (n_4192));
  NO2I1X1 g89337(.B (n_4133), .AN (\rs1_data[15]_39556 ), .Q (n_4190));
  NO2X1 g89338(.A (n_4137), .B (n_2423), .Q (n_4189));
  NO2X1 g89339(.A (n_4153), .B (n_2303), .Q (n_4188));
  NA2X1 g89340(.A (n_4137), .B (n_2423), .Q (n_4187));
  NO2X1 g89341(.A (n_4148), .B (n_6149), .Q (n_4186));
  NO2X1 g89342(.A (n_4143), .B (n_8366), .Q (n_4185));
  NO2I1X1 g89347(.B (n_4151), .AN (\rs1_data[30]_39526 ), .Q (n_4208));
  NA2X1 g89348(.A (n_4143), .B (n_8366), .Q (n_4207));
  NO2X1 g89349(.A (n_4153), .B (n_6141), .Q (n_4206));
  NA2X1 g89350(.A (n_4133), .B (n_2435), .Q (n_4205));
  NA2X1 g89351(.A (n_4134), .B (n_6127), .Q (n_4204));
  NO2X1 g89354(.A (n_4149), .B (n_2420), .Q (n_4203));
  NO2I1X1 g89355(.B (n_4150), .AN (n_6136), .Q (n_4202));
  NO2I1X1 g89357(.B (n_4152), .AN (\rs1_data[29]_39416 ), .Q (n_4201));
  NA2X1 g89359(.A (n_4149), .B (n_2420), .Q (n_4200));
  INX1 g89361(.A (n_4180), .Q (n_4181));
  INX1 g89365(.A (n_4171), .Q (n_4172));
  NA3X1 g89368(.A (n_4096), .B (n_2919), .C (n_2970), .Q (n_4169));
  NA2I1X1 g89370(.B (n_4119), .AN (\rs1_data[1]_39396 ), .Q (n_4167));
  NO2X1 g89371(.A (n_4146), .B (n_6132), .Q (n_4166));
  NA2I1X1 g89372(.B (n_4140), .AN (\rs1_data[24]_39336 ), .Q (n_4165));
  NO2X2 g89373(.A (n_2362), .B (n_2428), .Q (n_4164));
  NO2X1 g89376(.A (n_4134), .B (n_6127), .Q (n_4162));
  NA2I1X1 g89377(.B (n_8619), .AN (\rs1_data[26]_39356 ), .Q (n_4161));
  NA2I1X1 g89379(.B (n_4126), .AN (\rs1_data[12]_39516 ), .Q (n_4159));
  NO2I1X1 g89384(.B (n_4129), .AN (\rs1_data[23]_39326 ), .Q (n_4156));
  NO2X1 g89385(.A (n_4125), .B (n_2426), .Q (n_4155));
  NA2X2 g89387(.A (n_4125), .B (n_2426), .Q (n_4182));
  NA2X2 g89389(.A (n_4129), .B (n_2432), .Q (n_4180));
  NA2X2 g89390(.A (n_4128), .B (n_2429), .Q (n_2376));
  NA2X1 g89391(.A (n_4145), .B (n_501), .Q (n_4179));
  NO2I1X1 g89392(.B (n_4140), .AN (\rs1_data[24]_39336 ), .Q (n_4178));
  NO2X1 g89393(.A (n_4141), .B (\rs1_data[19]_39596 ), .Q (n_4177));
  NO2I1X1 g89394(.B (n_4145), .AN (\rs1_data[25]_39346 ), .Q (n_4176));
  NA2X1 g89395(.A (n_2365), .B (\rs1_data[3]_39426 ), .Q (n_4175));
  NO2I1X1 g89396(.B (n_4147), .AN (n_6132), .Q (n_4174));
  NA2X1 g89398(.A (n_8501), .B (n_2433), .Q (n_4173));
  NO2X2 g89399(.A (n_2369), .B (\rs1_data[21]_39616 ), .Q (n_4171));
  NO2I1X4 g89402(.B (n_4126), .AN (\rs1_data[12]_39516 ), .Q (n_4170));
  INX1 g89403(.A (n_4153), .Q (n_4154));
  INX1 g89405(.A (n_4147), .Q (n_4146));
  INX1 g89406(.A (n_4143), .Q (n_4144));
  INX1 g89407(.A (n_4142), .Q (n_4141));
  INX1 g89414(.A (n_4134), .Q (n_4135));
  INX1 g89416(.A (n_4131), .Q (n_4130));
  NO2X2 g89417(.A (n_4102), .B (n_4078), .Q (n_4153));
  NA3I1X4 g89418(.B (n_4089), .C (n_4091), .AN (n_4053), .Q (n_4152));
  NA3I1X2 g89419(.B (n_4087), .C (n_4092), .AN (n_4055), .Q (n_4151));
  NA3X2 g89420(.A (n_4088), .B (n_4083), .C (n_4049), .Q (n_4150));
  NA3I1X2 g89421(.B (n_4085), .C (n_4082), .AN (n_4046), .Q (n_4149));
  NO2X2 g89422(.A (n_4108), .B (n_4075), .Q (n_4148));
  NA3I1X4 g89423(.B (n_4073), .C (n_4066), .AN (n_4039), .Q (n_4147));
  NA3I1X4 g89424(.B (n_4072), .C (n_4065), .AN (n_4038), .Q (n_4145));
  NO2X2 g89425(.A (n_4107), .B (n_4093), .Q (n_4143));
  NA3X4 g89426(.A (n_4074), .B (n_4067), .C (n_4040), .Q (n_4142));
  NA3I1X4 g89427(.B (n_4071), .C (n_4064), .AN (n_4036), .Q (n_4140));
  NO2X4 g89429(.A (n_8700), .B (n_4079), .Q (n_2369));
  NA2X4 g89430(.A (n_4104), .B (n_4077), .Q (n_2368));
  NA3X4 g89431(.A (n_8505), .B (n_4084), .C (n_4048), .Q (n_4138));
  NA2X4 g89432(.A (n_4112), .B (n_4090), .Q (n_4137));
  NO2X4 g89433(.A (n_4109), .B (n_4080), .Q (n_4134));
  NA2X2 g89434(.A (n_4111), .B (n_4052), .Q (n_4133));
  NA2X4 g89435(.A (n_8502), .B (n_4094), .Q (n_4132));
  NO2X4 g89436(.A (n_4103), .B (n_4076), .Q (n_4131));
  INX3 g89437(.A (n_4124), .Q (n_4123));
  INX1 g89439(.A (n_2367), .Q (n_4121));
  INX1 g89444(.A (n_8501), .Q (n_4116));
  INX1 g89445(.A (n_2364), .Q (n_4115));
  BUX1 g89447(.A (n_2363), .Q (n_2364));
  INX1 g89449(.A (n_2362), .Q (n_4114));
  ON21X1 g89452(.A (n_4050), .B (n_3085), .C (n_2503), .Q (n_8191));
  ON21X1 g89453(.A (n_4051), .B (n_3086), .C (n_2503), .Q (n_8183));
  ON21X1 g89454(.A (n_4051), .B (n_3084), .C (n_2503), .Q (n_8187));
  ON21X1 g89455(.A (n_4051), .B (n_3085), .C (n_2503), .Q (n_8188));
  ON21X1 g89456(.A (n_4050), .B (n_3086), .C (n_2503), .Q (n_8180));
  ON21X1 g89457(.A (n_4050), .B (n_3087), .C (n_2503), .Q (n_8196));
  ON21X1 g89458(.A (n_4051), .B (n_3087), .C (n_2503), .Q (n_8198));
  ON21X1 g89459(.A (n_4050), .B (n_3084), .C (n_2503), .Q (n_8202));
  NA3X4 g89460(.A (n_4070), .B (n_4059), .C (n_4026), .Q (n_4129));
  NA2X4 g89461(.A (n_4100), .B (n_4056), .Q (n_4128));
  NA2X4 g89462(.A (n_8504), .B (n_4063), .Q (n_4127));
  NA3X2 g89463(.A (n_4044), .B (n_4033), .C (n_4016), .Q (n_4126));
  NA3X2 g89464(.A (n_4062), .B (n_4035), .C (n_4019), .Q (n_4125));
  NA2X4 g89465(.A (n_4101), .B (n_4045), .Q (n_4124));
  NA3X4 g89466(.A (n_4097), .B (n_4014), .C (n_4011), .Q (n_2367));
  NA3X4 g89467(.A (n_4023), .B (n_4015), .C (n_4009), .Q (n_4119));
  NA3X4 g89468(.A (n_4025), .B (n_4013), .C (n_4010), .Q (n_4118));
  NA3X2 g89470(.A (n_4069), .B (n_4043), .C (n_4022), .Q (n_2363));
  NA3X4 g89471(.A (n_4068), .B (n_4042), .C (n_4021), .Q (n_2362));
  NO3X1 g89472(.A (n_4054), .B (n_3980), .C (n_3984), .Q (n_4112));
  NO3X2 g89473(.A (n_4095), .B (n_3979), .C (n_3983), .Q (n_4111));
  NA3X1 g89475(.A (n_4031), .B (n_8514), .C (n_8512), .Q (n_4109));
  NA3X1 g89476(.A (n_4041), .B (n_8515), .C (n_8513), .Q (n_4108));
  NA3X1 g89477(.A (n_4037), .B (n_2361), .C (n_8678), .Q (n_4107));
  NO2X2 g89480(.A (n_4061), .B (n_4032), .Q (n_4104));
  NA2X1 g89481(.A (n_4057), .B (n_4028), .Q (n_4103));
  NA3X1 g89482(.A (n_4027), .B (n_2359), .C (n_2360), .Q (n_4102));
  NO3X4 g89483(.A (n_4017), .B (n_3916), .C (n_8516), .Q (n_4101));
  NO2X2 g89484(.A (n_8506), .B (n_4018), .Q (n_4100));
  ON21X1 g89486(.A (n_3947), .B (n_3078), .C (n_2503), .Q (n_8201));
  ON21X1 g89487(.A (n_3945), .B (n_3078), .C (n_2503), .Q (n_8199));
  ON21X1 g89488(.A (n_3946), .B (n_3083), .C (n_2503), .Q (n_8197));
  ON21X1 g89489(.A (n_3947), .B (n_3083), .C (n_2503), .Q (n_8194));
  ON21X1 g89490(.A (n_3945), .B (n_3083), .C (n_2503), .Q (n_8190));
  ON21X1 g89491(.A (n_3946), .B (n_3077), .C (n_2503), .Q (n_8185));
  ON21X1 g89492(.A (n_3947), .B (n_3077), .C (n_2503), .Q (n_8182));
  ON21X1 g89493(.A (n_3945), .B (n_3077), .C (n_2503), .Q (n_8181));
  ON21X1 g89494(.A (n_3946), .B (n_3079), .C (n_2503), .Q (n_8178));
  ON21X1 g89495(.A (n_3947), .B (n_3079), .C (n_2503), .Q (n_8175));
  ON21X1 g89496(.A (n_3945), .B (n_3079), .C (n_2503), .Q (n_8174));
  ON21X1 g89497(.A (n_3946), .B (n_3078), .C (n_2503), .Q (n_8171));
  ON21X1 g89499(.A (n_3948), .B (n_3083), .C (n_2503), .Q (n_8186));
  ON21X1 g89500(.A (n_3948), .B (n_3077), .C (n_2503), .Q (n_8179));
  ON21X1 g89501(.A (n_3948), .B (n_3079), .C (n_2503), .Q (n_8172));
  NO3X2 g89502(.A (n_3898), .B (n_3660), .C (n_3882), .Q (n_4097));
  ON21X0 g89503(.A (n_3943), .B (n_3180), .C (n_2503), .Q (n_8203));
  ON21X1 g89504(.A (n_3944), .B (n_3180), .C (n_2503), .Q (n_8200));
  ON21X0 g89505(.A (n_3943), .B (n_3184), .C (n_2503), .Q (n_8195));
  ON21X1 g89506(.A (n_3944), .B (n_3184), .C (n_2503), .Q (n_8193));
  ON21X0 g89507(.A (n_3943), .B (n_3183), .C (n_2503), .Q (n_8192));
  ON21X1 g89508(.A (n_3944), .B (n_3183), .C (n_2503), .Q (n_8189));
  ON21X0 g89509(.A (n_3943), .B (n_3181), .C (n_2503), .Q (n_8176));
  ON21X1 g89510(.A (n_3944), .B (n_3181), .C (n_2503), .Q (n_8173));
  AN31X1 g89511(.A (n_2487), .B (n_2609), .C (n_2764), .D (n_4007), .Q
       (n_4096));
  NA3X1 g89512(.A (n_3921), .B (n_3735), .C (n_3736), .Q (n_4095));
  NO2X1 g89513(.A (n_3999), .B (n_3989), .Q (n_4094));
  NA3X1 g89514(.A (n_3966), .B (n_2349), .C (n_2348), .Q (n_4093));
  AND4X1 g89515(.A (n_3810), .B (n_3797), .C (n_3811), .D (n_3798), .Q
       (n_4092));
  AND4X1 g89516(.A (n_3806), .B (n_3793), .C (n_3807), .D (n_3794), .Q
       (n_4091));
  AND6X2 g89517(.A (n_8530), .B (n_3773), .C (n_3494), .D (n_3473), .E
       (n_3487), .F (n_3466), .Q (n_4090));
  NO2X1 g89518(.A (n_8509), .B (n_3988), .Q (n_4089));
  NO2X1 g89519(.A (n_8510), .B (n_3987), .Q (n_4088));
  NO3X1 g89520(.A (n_3986), .B (n_3854), .C (n_3856), .Q (n_4087));
  NO3X1 g89522(.A (n_3977), .B (n_3858), .C (n_3853), .Q (n_4085));
  NO2X1 g89523(.A (n_3978), .B (n_3976), .Q (n_4084));
  AND4X1 g89524(.A (n_3800), .B (n_3788), .C (n_3801), .D (n_3779), .Q
       (n_4083));
  AND4X1 g89525(.A (n_3814), .B (n_3786), .C (n_3815), .D (n_3787), .Q
       (n_4082));
  NA3X2 g89527(.A (n_3955), .B (n_2347), .C (n_8534), .Q (n_4080));
  NA3X2 g89528(.A (n_3954), .B (n_3839), .C (n_3836), .Q (n_4079));
  NA3X2 g89529(.A (n_3953), .B (n_2353), .C (n_2351), .Q (n_4078));
  NO2X2 g89530(.A (n_3994), .B (n_3952), .Q (n_4077));
  NA3X2 g89531(.A (n_3951), .B (n_2352), .C (n_3835), .Q (n_4076));
  NA2X2 g89532(.A (n_3993), .B (n_3965), .Q (n_4075));
  NO2X2 g89533(.A (n_3995), .B (n_3964), .Q (n_4074));
  NO3X1 g89534(.A (n_3963), .B (n_3842), .C (n_3845), .Q (n_4073));
  NO2X2 g89535(.A (n_3992), .B (n_3962), .Q (n_4072));
  NO2X2 g89536(.A (n_8511), .B (n_3961), .Q (n_4071));
  NO3X2 g89537(.A (n_3950), .B (n_3834), .C (n_3838), .Q (n_4070));
  NO3X2 g89538(.A (n_3932), .B (n_3831), .C (n_3833), .Q (n_4069));
  NO3X2 g89539(.A (n_3933), .B (n_3830), .C (n_3832), .Q (n_4068));
  NO2X1 g89540(.A (n_3973), .B (n_3968), .Q (n_4067));
  NO2X1 g89541(.A (n_3972), .B (n_3958), .Q (n_4066));
  NO2X1 g89542(.A (n_3971), .B (n_3957), .Q (n_4065));
  NO2X1 g89543(.A (n_3969), .B (n_3967), .Q (n_4064));
  NO3X2 g89544(.A (n_3925), .B (n_3824), .C (n_3829), .Q (n_4063));
  NO3X1 g89545(.A (n_3926), .B (n_3817), .C (n_3818), .Q (n_4062));
  NA3X1 g89546(.A (n_8508), .B (n_3615), .C (n_3710), .Q (n_4061));
  NO2X1 g89548(.A (n_3938), .B (n_3934), .Q (n_4059));
  NA3X1 g89549(.A (n_3940), .B (n_3704), .C (n_3707), .Q (n_4058));
  NO2X1 g89550(.A (n_3939), .B (n_3935), .Q (n_4057));
  AND6X2 g89551(.A (n_8535), .B (n_3588), .C (n_3353), .D (n_3324), .E
       (n_3329), .F (n_3354), .Q (n_4056));
  NA3X1 g89552(.A (n_3924), .B (n_3740), .C (n_3741), .Q (n_4055));
  NA3X1 g89553(.A (n_3923), .B (n_3738), .C (n_3739), .Q (n_4054));
  NA3X1 g89554(.A (n_3922), .B (n_3742), .C (n_3737), .Q (n_4053));
  NO3X1 g89555(.A (n_3990), .B (n_3851), .C (n_3852), .Q (n_4052));
  AND3X1 g89556(.A (n_3920), .B (n_3731), .C (n_3732), .Q (n_4049));
  AND4X1 g89557(.A (n_3713), .B (n_3733), .C (n_3734), .D (n_3632), .Q
       (n_4048));
  NA3X1 g89559(.A (n_3928), .B (n_3777), .C (n_3778), .Q (n_4046));
  NO3X4 g89560(.A (n_3931), .B (n_3823), .C (n_3828), .Q (n_4045));
  NO3X2 g89561(.A (n_3930), .B (n_3822), .C (n_3827), .Q (n_4044));
  AND4X1 g89562(.A (n_3642), .B (n_3646), .C (n_3643), .D (n_3647), .Q
       (n_4043));
  NO2X1 g89563(.A (n_3929), .B (n_3927), .Q (n_4042));
  AND4X1 g89564(.A (n_3727), .B (n_3728), .C (n_3655), .D (n_3584), .Q
       (n_4041));
  NO2X1 g89565(.A (n_3949), .B (n_3907), .Q (n_4040));
  NA3X1 g89566(.A (n_8517), .B (n_3723), .C (n_3724), .Q (n_4039));
  NA3X1 g89567(.A (n_3905), .B (n_3721), .C (n_3722), .Q (n_4038));
  AND4X1 g89568(.A (n_3719), .B (n_3720), .C (n_3653), .D (n_3582), .Q
       (n_4037));
  NA3X1 g89569(.A (n_8518), .B (n_3717), .C (n_3718), .Q (n_4036));
  NO2X1 g89570(.A (n_3918), .B (n_3913), .Q (n_4035));
  NO2X1 g89572(.A (n_3915), .B (n_3910), .Q (n_4033));
  NA3X1 g89573(.A (n_8519), .B (n_3682), .C (n_3683), .Q (n_4032));
  AND4X1 g89574(.A (n_3680), .B (n_3681), .C (n_3639), .D (n_3572), .Q
       (n_4031));
  NA3X1 g89575(.A (n_3902), .B (n_3675), .C (n_3678), .Q (n_4030));
  NO2X1 g89577(.A (n_3937), .B (n_3900), .Q (n_4028));
  AND4X1 g89578(.A (n_3666), .B (n_3667), .C (n_3628), .D (n_3574), .Q
       (n_4027));
  AND4X1 g89579(.A (n_3663), .B (n_3664), .C (n_3636), .D (n_3570), .Q
       (n_4026));
  NO3X2 g89580(.A (n_3899), .B (n_3661), .C (n_3652), .Q (n_4025));
  NO2X2 g89581(.A (n_3908), .B (n_3897), .Q (n_4024));
  NO2X2 g89582(.A (n_3909), .B (n_8621), .Q (n_4023));
  AND4X1 g89583(.A (n_3603), .B (n_3604), .C (n_3567), .D (n_3556), .Q
       (n_4022));
  AND4X1 g89584(.A (n_3601), .B (n_3602), .C (n_3566), .D (n_3555), .Q
       (n_4021));
  AND4X1 g89586(.A (n_3599), .B (n_3598), .C (n_3565), .D (n_3542), .Q
       (n_4019));
  NA3X1 g89587(.A (n_2357), .B (n_3596), .C (n_3597), .Q (n_4018));
  NA3X2 g89588(.A (n_3894), .B (n_8556), .C (n_3593), .Q (n_4017));
  AND4X1 g89589(.A (n_3591), .B (n_3590), .C (n_3561), .D (n_3538), .Q
       (n_4016));
  NO3X2 g89590(.A (n_3891), .B (n_3558), .C (n_3545), .Q (n_4015));
  NO3X2 g89591(.A (n_3893), .B (n_3560), .C (n_3553), .Q (n_4014));
  NO3X2 g89592(.A (n_3892), .B (n_3549), .C (n_3550), .Q (n_4013));
  NO3X2 g89594(.A (n_3886), .B (n_3267), .C (n_3530), .Q (n_4011));
  NO2X2 g89595(.A (n_3888), .B (n_3883), .Q (n_4010));
  NO2X2 g89596(.A (n_3887), .B (n_3884), .Q (n_4009));
  NA3X1 g89597(.A (n_8522), .B (n_3532), .C (n_3535), .Q (n_4008));
  NO3I1X1 g89598(.B (n_8523), .C (n_8157), .AN (system_type), .Q
       (n_4007));
  OR2X1 g89599(.A (n_3943), .B (n_2804), .Q (n_4051));
  NA2X1 g89600(.A (n_2282), .B (n_2805), .Q (n_4050));
  INX6 g89601(.A (n_8655), .Q (n_7383));
  INX4 g89602(.A (inc_ADD_UNS_OP5491_6_n_2669), .Q (n_7381));
  INX4 g89603(.A (n_8657), .Q (n_7395));
  INX3 g89606(.A (n_4002), .Q (n_7387));
  INX3 g89607(.A (n_4001), .Q (n_7386));
  INX3 g89608(.A (n_4000), .Q (n_7388));
  NA2X2 g89611(.A (n_3874), .B (n_2669), .Q (n_7379));
  NA2X2 g89613(.A (n_3877), .B (n_2670), .Q (n_7635));
  NA2X2 g89614(.A (n_3875), .B (n_2664), .Q (n_7378));
  NA2X4 g89615(.A (n_3873), .B (n_2666), .Q (n_7380));
  NA2X2 g89616(.A (n_3872), .B (n_2667), .Q (n_7384));
  OA22X4 g89617(.A (n_2660), .B (n_2346), .C (n_501), .D (n_2588), .Q
       (inc_ADD_UNS_OP5491_6_n_2669));
  NA2X4 g89619(.A (n_3871), .B (n_2671), .Q (n_7376));
  NO2X4 g89622(.A (n_3866), .B (n_2661), .Q (n_4002));
  NO2X2 g89623(.A (n_8527), .B (n_2320), .Q (n_4001));
  NO2X2 g89624(.A (n_8528), .B (n_2319), .Q (n_4000));
  NA2X2 g89625(.A (n_3864), .B (n_2658), .Q (n_7399));
  NA2X4 g89626(.A (n_3860), .B (n_8567), .Q (n_8208));
  NA2X4 g89628(.A (n_3859), .B (n_2650), .Q (n_7389));
  NA3X1 g89629(.A (n_8529), .B (n_3470), .C (n_3455), .Q (n_3999));
  NA3X2 g89632(.A (n_3846), .B (n_3442), .C (n_3512), .Q (n_3996));
  NA3X2 g89633(.A (n_8532), .B (n_3429), .C (n_3453), .Q (n_3995));
  NA3X1 g89634(.A (n_8533), .B (n_3444), .C (n_3401), .Q (n_3994));
  AND4X1 g89635(.A (n_3454), .B (n_3431), .C (n_3432), .D (n_3419), .Q
       (n_3993));
  NA3X1 g89636(.A (n_8531), .B (n_3451), .C (n_3426), .Q (n_3992));
  NA3X2 g89638(.A (n_8538), .B (n_3463), .C (n_3409), .Q (n_3990));
  NA3X1 g89639(.A (n_3781), .B (n_3456), .C (n_3496), .Q (n_3989));
  NA3X1 g89640(.A (n_8539), .B (n_3465), .C (n_3436), .Q (n_3988));
  NA3X1 g89641(.A (n_8540), .B (n_3462), .C (n_3435), .Q (n_3987));
  NA3X1 g89642(.A (n_8541), .B (n_3457), .C (n_3433), .Q (n_3986));
  NA2X1 g89644(.A (n_3795), .B (n_3796), .Q (n_3984));
  NA2X1 g89645(.A (n_3791), .B (n_3792), .Q (n_3983));
  NA2X1 g89646(.A (n_3799), .B (n_3790), .Q (n_3982));
  NA2X1 g89647(.A (n_3812), .B (n_3813), .Q (n_3981));
  NA2X1 g89648(.A (n_3808), .B (n_3809), .Q (n_3980));
  NA2X1 g89649(.A (n_3804), .B (n_3805), .Q (n_3979));
  NA2X1 g89650(.A (n_3802), .B (n_3881), .Q (n_3978));
  NA3X1 g89651(.A (n_8536), .B (n_3477), .C (n_3469), .Q (n_3977));
  NA2X1 g89652(.A (n_3789), .B (n_3780), .Q (n_3976));
  NA2X1 g89655(.A (n_3760), .B (n_3761), .Q (n_3973));
  NA2X1 g89656(.A (n_3758), .B (n_3759), .Q (n_3972));
  NA2X1 g89657(.A (n_3756), .B (n_3757), .Q (n_3971));
  NA2X1 g89659(.A (n_3752), .B (n_3753), .Q (n_3969));
  NA2X1 g89660(.A (n_3748), .B (n_8543), .Q (n_3968));
  NA2X1 g89661(.A (n_3743), .B (n_3744), .Q (n_3967));
  NO2X1 g89662(.A (n_3825), .B (n_8542), .Q (n_3966));
  NO2X1 g89663(.A (n_3826), .B (n_8545), .Q (n_3965));
  NA3X1 g89664(.A (n_8546), .B (n_3399), .C (n_3418), .Q (n_3964));
  NA3X2 g89665(.A (n_8547), .B (n_3398), .C (n_3416), .Q (n_3963));
  NA3X1 g89666(.A (n_3669), .B (n_3397), .C (n_3414), .Q (n_3962));
  NA3X2 g89667(.A (n_8701), .B (n_3395), .C (n_3411), .Q (n_3961));
  NA2X1 g89670(.A (n_3747), .B (n_3768), .Q (n_3958));
  NA2X1 g89671(.A (n_3746), .B (n_3767), .Q (n_3957));
  NA3X1 g89673(.A (n_3685), .B (n_3378), .C (n_3500), .Q (n_3956));
  NO2X1 g89674(.A (n_3821), .B (n_8544), .Q (n_3955));
  NO2X1 g89675(.A (n_3820), .B (n_3679), .Q (n_3954));
  NO2X1 g89676(.A (n_3819), .B (n_8548), .Q (n_3953));
  NA3X1 g89677(.A (n_3373), .B (n_3662), .C (n_3509), .Q (n_3952));
  NO2X1 g89678(.A (n_3816), .B (n_8537), .Q (n_3951));
  NA3X2 g89679(.A (n_8551), .B (n_3374), .C (n_3507), .Q (n_3950));
  NA2X1 g89680(.A (n_3725), .B (n_3726), .Q (n_3949));
  NA2X4 g89681(.A (n_3876), .B (n_2668), .Q (n_7377));
  INX1 g89682(.A (n_2282), .Q (n_3944));
  NA2X1 g89683(.A (n_3676), .B (n_3677), .Q (n_3942));
  NA2X1 g89684(.A (n_3694), .B (n_3695), .Q (n_3941));
  NO2X1 g89685(.A (n_3692), .B (n_3693), .Q (n_3940));
  NA2X1 g89686(.A (n_3690), .B (n_3691), .Q (n_3939));
  NA2X1 g89688(.A (n_3686), .B (n_3687), .Q (n_3938));
  NA2X1 g89689(.A (n_3670), .B (n_3671), .Q (n_3937));
  NA2X1 g89690(.A (n_3705), .B (n_3706), .Q (n_3936));
  NA2X1 g89691(.A (n_3702), .B (n_3703), .Q (n_3935));
  NA2X1 g89693(.A (n_3698), .B (n_3699), .Q (n_3934));
  NA3X1 g89694(.A (n_3708), .B (n_3346), .C (n_3315), .Q (n_3933));
  NA3X1 g89695(.A (n_3600), .B (n_3362), .C (n_3287), .Q (n_3932));
  NA3X2 g89696(.A (n_8680), .B (n_3317), .C (n_3276), .Q (n_3931));
  NA3X1 g89697(.A (n_8681), .B (n_3316), .C (n_3275), .Q (n_3930));
  NA2X1 g89698(.A (n_3640), .B (n_3641), .Q (n_3929));
  NO3X1 g89699(.A (n_3648), .B (n_3344), .C (n_3345), .Q (n_3928));
  NA2X1 g89700(.A (n_8553), .B (n_8552), .Q (n_3927));
  NA3X1 g89701(.A (n_3589), .B (n_3311), .C (n_3356), .Q (n_3926));
  NA3X1 g89702(.A (n_3587), .B (n_3318), .C (n_3310), .Q (n_3925));
  NO2X1 g89703(.A (n_3716), .B (n_3635), .Q (n_3924));
  NO2X1 g89704(.A (n_3715), .B (n_3634), .Q (n_3923));
  NO2X1 g89705(.A (n_3714), .B (n_3633), .Q (n_3922));
  AND3X1 g89706(.A (n_8554), .B (n_3312), .C (n_3313), .Q (n_3921));
  NO2X1 g89707(.A (n_3712), .B (n_3626), .Q (n_3920));
  NA2X1 g89709(.A (n_3613), .B (n_3614), .Q (n_3918));
  NA2X1 g89711(.A (n_3609), .B (n_3610), .Q (n_3917));
  NA2X1 g89712(.A (n_3608), .B (n_3607), .Q (n_3916));
  NA2X1 g89713(.A (n_3605), .B (n_3606), .Q (n_3915));
  NA2X1 g89715(.A (n_3624), .B (n_3625), .Q (n_3913));
  NO2X1 g89716(.A (n_3622), .B (n_3623), .Q (n_3912));
  NA2X1 g89717(.A (n_3620), .B (n_3621), .Q (n_3911));
  NA2X1 g89718(.A (n_3616), .B (n_3617), .Q (n_3910));
  NA3X1 g89719(.A (n_8550), .B (n_3263), .C (n_3260), .Q (n_3909));
  NA3X1 g89720(.A (n_3651), .B (n_3261), .C (n_3262), .Q (n_3908));
  NA2X1 g89721(.A (n_3658), .B (n_3581), .Q (n_3907));
  NO2X1 g89723(.A (n_3657), .B (n_3579), .Q (n_3905));
  NO2X2 g89726(.A (n_3638), .B (n_3573), .Q (n_3902));
  NA2X1 g89728(.A (n_3629), .B (n_8558), .Q (n_3900));
  NA3X2 g89729(.A (n_8557), .B (n_3255), .C (n_3270), .Q (n_3899));
  NA3X1 g89730(.A (n_3578), .B (n_3271), .C (n_3233), .Q (n_3898));
  NA3X2 g89731(.A (n_3268), .B (n_8682), .C (n_3240), .Q (n_3897));
  NO2X2 g89735(.A (n_3562), .B (n_3539), .Q (n_3894));
  NA2X1 g89736(.A (n_3551), .B (n_3552), .Q (n_3893));
  NA2X1 g89737(.A (n_3547), .B (n_3548), .Q (n_3892));
  NA2X1 g89738(.A (n_3559), .B (n_3546), .Q (n_3891));
  NA2X1 g89741(.A (n_3537), .B (n_3534), .Q (n_3888));
  NA2X1 g89742(.A (n_3533), .B (n_3536), .Q (n_3887));
  NA2X1 g89743(.A (n_3528), .B (n_3529), .Q (n_3886));
  NO3I1X1 g89744(.B (n_8300), .C (n_2586), .AN (n_7371), .Q (n_7861));
  NA2X1 g89746(.A (n_3526), .B (n_3524), .Q (n_3884));
  NA2X1 g89747(.A (n_3527), .B (n_3523), .Q (n_3883));
  NA2X1 g89748(.A (n_3531), .B (n_3234), .Q (n_3882));
  NA3X1 g89750(.A (n_3709), .B (n_2504), .C (n_2417), .Q (n_3948));
  NA3X1 g89751(.A (n_3709), .B (n_2602), .C (n_2417), .Q (n_3947));
  NA3X1 g89752(.A (n_3709), .B (n_2602), .C (\instruction[7]_39642 ),
       .Q (n_3946));
  NA3X1 g89753(.A (n_3709), .B (n_2504), .C (\instruction[7]_39642 ),
       .Q (n_3945));
  NA3X1 g89755(.A (n_3006), .B (n_3179), .C (\instruction[7]_39642 ),
       .Q (n_3943));
  INX4 g89756(.A (n_3880), .Q (n_7391));
  INX3 g89757(.A (inc_ADD_UNS_OP_5_n_3766), .Q (n_7392));
  INX4 g89758(.A (inc_ADD_UNS_OP5491_6_n_2675), .Q (n_7393));
  INX8 g89760(.A (n_3863), .Q (n_7632));
  INX6 g89761(.A (n_3862), .Q (n_7398));
  AN22X1 g89763(.A (n_3165), .B (n_6956), .C (n_3173), .D (n_6954), .Q
       (n_3881));
  OA21X4 g89764(.A (n_2435), .B (n_2588), .C (n_3522), .Q (n_3880));
  OA21X4 g89765(.A (n_2425), .B (n_2588), .C (n_3521), .Q
       (inc_ADD_UNS_OP_5_n_3766));
  AND2X4 g89766(.A (n_3520), .B (n_2662), .Q
       (inc_ADD_UNS_OP5491_6_n_2675));
  NA2X2 g89767(.A (n_3519), .B (n_2656), .Q (n_7394));
  NA2X2 g89768(.A (n_3518), .B (n_2659), .Q (n_7400));
  ON21X1 g89770(.A (n_2543), .B (n_2590), .C (csr_data_out[31]), .Q
       (n_3877));
  ON21X1 g89771(.A (n_2539), .B (n_2590), .C (csr_data_out[29]), .Q
       (n_3876));
  ON21X1 g89772(.A (n_2545), .B (n_2590), .C (csr_data_out[28]), .Q
       (n_3875));
  ON21X1 g89773(.A (n_2541), .B (n_2590), .C (csr_data_out[27]), .Q
       (n_3874));
  ON21X1 g89774(.A (n_2544), .B (n_2590), .C (csr_data_out[26]), .Q
       (n_3873));
  ON21X1 g89775(.A (n_2540), .B (n_2590), .C (csr_data_out[22]), .Q
       (n_3872));
  ON21X1 g89776(.A (n_2538), .B (n_2590), .C (csr_data_out[30]), .Q
       (n_3871));
  NO2I1X2 g89781(.B (n_2676), .AN (csr_data_out[19]), .Q (n_3866));
  ON21X1 g89783(.A (n_2531), .B (n_2590), .C (csr_data_out[7]), .Q
       (n_3864));
  NO2X4 g89785(.A (n_3515), .B (n_2713), .Q (n_3863));
  NO2X4 g89786(.A (n_3517), .B (n_2318), .Q (n_3862));
  NA2X4 g89787(.A (n_3513), .B (n_2649), .Q (n_7401));
  NA2X4 g89788(.A (n_3514), .B (n_2648), .Q (n_7397));
  ON31X1 g89790(.A (n_2507), .B (n_2582), .C (n_2584), .D
       (csr_data_out[3]), .Q (n_3860));
  ON21X1 g89791(.A (n_2523), .B (n_2590), .C (csr_data_out[17]), .Q
       (n_3859));
  NA2X1 g89792(.A (n_3479), .B (n_3478), .Q (n_3858));
  AND2X2 g89794(.A (n_3493), .B (n_3464), .Q (n_3857));
  NA2X1 g89795(.A (n_3489), .B (n_3474), .Q (n_3856));
  NA2X1 g89797(.A (n_3483), .B (n_3458), .Q (n_3855));
  NA2X1 g89798(.A (n_3482), .B (n_3468), .Q (n_3854));
  NA2X1 g89799(.A (n_3495), .B (n_3480), .Q (n_3853));
  NA2X1 g89800(.A (n_3461), .B (n_3472), .Q (n_3852));
  NA2X1 g89801(.A (n_3485), .B (n_3492), .Q (n_3851));
  NO2X1 g89802(.A (n_3484), .B (n_3491), .Q (n_3850));
  NA2X1 g89804(.A (n_3490), .B (n_3471), .Q (n_3848));
  NO2X1 g89808(.A (n_3406), .B (n_3501), .Q (n_3846));
  NA2X1 g89809(.A (n_3427), .B (n_3415), .Q (n_3845));
  NA2X1 g89814(.A (n_3452), .B (n_3428), .Q (n_3842));
  NO2X1 g89816(.A (n_3449), .B (n_3422), .Q (n_3841));
  AND2X1 g89820(.A (n_3306), .B (n_3503), .Q (n_3839));
  NA2X1 g89821(.A (n_3381), .B (n_3508), .Q (n_3838));
  NO2X1 g89823(.A (n_3441), .B (n_3404), .Q (n_3836));
  AND2X1 g89824(.A (n_3439), .B (n_3403), .Q (n_3835));
  NA2X1 g89825(.A (n_3438), .B (n_3402), .Q (n_3834));
  NA2X1 g89826(.A (n_3360), .B (n_3367), .Q (n_3833));
  NA2X1 g89827(.A (n_3359), .B (n_3365), .Q (n_3832));
  NA2X1 g89828(.A (n_3358), .B (n_3366), .Q (n_3831));
  NA2X1 g89829(.A (n_3357), .B (n_3364), .Q (n_3830));
  NA2X1 g89830(.A (n_3328), .B (n_3352), .Q (n_3829));
  NA2X1 g89831(.A (n_3350), .B (n_3327), .Q (n_3828));
  NA2X1 g89832(.A (n_3326), .B (n_3348), .Q (n_3827));
  NA2X1 g89833(.A (n_3420), .B (n_3400), .Q (n_3826));
  NA2X1 g89834(.A (n_3412), .B (n_3396), .Q (n_3825));
  NA2X1 g89835(.A (n_3323), .B (n_3351), .Q (n_3824));
  NA2X1 g89836(.A (n_3322), .B (n_3349), .Q (n_3823));
  NA2X1 g89837(.A (n_3321), .B (n_3347), .Q (n_3822));
  NA2X1 g89838(.A (n_3379), .B (n_3498), .Q (n_3821));
  NA2X1 g89839(.A (n_3502), .B (n_8560), .Q (n_3820));
  NA2X1 g89840(.A (n_3375), .B (n_3505), .Q (n_3819));
  NA2X1 g89841(.A (n_3355), .B (n_3330), .Q (n_3818));
  NA2X1 g89842(.A (n_3320), .B (n_3325), .Q (n_3817));
  NA2X1 g89843(.A (n_3376), .B (n_3361), .Q (n_3816));
  AN22X1 g89844(.A (n_3171), .B (n_7237), .C (n_3173), .D (n_7233), .Q
       (n_3815));
  AN22X1 g89845(.A (n_3170), .B (n_7239), .C (n_3165), .D (n_7235), .Q
       (n_3814));
  AN21X1 g89846(.A (n_3171), .B (n_6927), .C (n_3387), .Q (n_3813));
  AN22X1 g89847(.A (n_3170), .B (n_6929), .C (n_3165), .D (n_6925), .Q
       (n_3812));
  AN22X1 g89848(.A (n_3171), .B (n_6896), .C (n_3165), .D (n_6894), .Q
       (n_3811));
  AN22X1 g89849(.A (n_3170), .B (n_6898), .C (n_3173), .D (n_6892), .Q
       (n_3810));
  AN22X1 g89850(.A (n_3171), .B (n_6400), .C (n_3165), .D (n_6398), .Q
       (n_3809));
  AN22X1 g89851(.A (n_3170), .B (n_6402), .C (n_3173), .D (n_6396), .Q
       (n_3808));
  AN22X1 g89852(.A (n_3171), .B (n_6555), .C (n_3165), .D (n_6553), .Q
       (n_3807));
  AN22X1 g89853(.A (n_3170), .B (n_6557), .C (n_3173), .D (n_6551), .Q
       (n_3806));
  AN21X1 g89854(.A (n_3171), .B (n_6989), .C (n_3386), .Q (n_3805));
  AN21X1 g89855(.A (n_3170), .B (n_6991), .C (n_3385), .Q (n_3804));
  AN22X1 g89857(.A (n_3170), .B (n_6960), .C (n_3171), .D (n_6958), .Q
       (n_3802));
  AN22X1 g89858(.A (n_3165), .B (n_6429), .C (n_3173), .D (n_6427), .Q
       (n_3801));
  AN22X1 g89859(.A (n_3170), .B (n_6433), .C (n_3171), .D (n_6431), .Q
       (n_3800));
  AN21X1 g89860(.A (n_3167), .B (n_6930), .C (n_3392), .Q (n_3799));
  AN22X1 g89861(.A (n_3177), .B (n_6897), .C (n_3175), .D (n_6895), .Q
       (n_3798));
  AN22X1 g89862(.A (n_3167), .B (n_6899), .C (n_2300), .D (n_6893), .Q
       (n_3797));
  AN22X1 g89863(.A (n_3177), .B (n_6401), .C (n_3175), .D (n_6399), .Q
       (n_3796));
  AN22X1 g89864(.A (n_3167), .B (n_6403), .C (n_2300), .D (n_6397), .Q
       (n_3795));
  AN22X1 g89865(.A (n_3177), .B (n_6556), .C (n_3175), .D (n_6554), .Q
       (n_3794));
  AN22X1 g89866(.A (n_3167), .B (n_6558), .C (n_2300), .D (n_6552), .Q
       (n_3793));
  NO2X1 g89867(.A (n_3390), .B (n_3391), .Q (n_3792));
  AN21X1 g89868(.A (n_3167), .B (n_6992), .C (n_3389), .Q (n_3791));
  AN21X1 g89869(.A (n_3177), .B (n_6928), .C (n_3393), .Q (n_3790));
  AN22X1 g89870(.A (n_3167), .B (n_6961), .C (n_3177), .D (n_6959), .Q
       (n_3789));
  AN22X1 g89871(.A (n_3167), .B (n_6434), .C (n_3177), .D (n_6432), .Q
       (n_3788));
  AN22X1 g89872(.A (n_3177), .B (n_7238), .C (n_2300), .D (n_7234), .Q
       (n_3787));
  AN22X1 g89873(.A (n_3167), .B (n_7240), .C (n_3175), .D (n_7236), .Q
       (n_3786));
  AN211X1 g89878(.A (n_3075), .B (n_6916), .C (n_3218), .D (n_3190), .Q
       (n_3781));
  AN21X1 g89879(.A (n_3175), .B (n_6957), .C (n_3388), .Q (n_3780));
  AN22X1 g89880(.A (n_3175), .B (n_6430), .C (n_2300), .D (n_6428), .Q
       (n_3779));
  AN22X1 g89881(.A (n_3154), .B (n_7245), .C (n_3152), .D (n_7243), .Q
       (n_3778));
  AN22X1 g89882(.A (n_3156), .B (n_7247), .C (n_3163), .D (n_7241), .Q
       (n_3777));
  AN221X1 g89886(.A (n_6388), .B (n_3073), .C (n_6389), .D (n_3075), .E
       (n_3149), .Q (n_3773));
  AO22X1 g89889(.A (n_3175), .B (n_6740), .C (n_2300), .D (n_6738), .Q
       (n_3770));
  AN22X1 g89891(.A (n_3175), .B (n_7019), .C (n_2300), .D (n_7017), .Q
       (n_3768));
  AN22X1 g89892(.A (n_3175), .B (n_6337), .C (n_2300), .D (n_6335), .Q
       (n_3767));
  AN22X1 g89893(.A (n_3175), .B (n_7050), .C (n_2300), .D (n_7048), .Q
       (n_3766));
  NA2X1 g89895(.A (n_3338), .B (n_3337), .Q (n_3764));
  NA2X1 g89896(.A (n_3335), .B (n_3336), .Q (n_3763));
  AN22X1 g89898(.A (n_3171), .B (n_7113), .C (n_3165), .D (n_7111), .Q
       (n_3761));
  AN22X1 g89899(.A (n_3170), .B (n_7115), .C (n_3173), .D (n_7109), .Q
       (n_3760));
  AN22X1 g89900(.A (n_3165), .B (n_7018), .C (n_3173), .D (n_7016), .Q
       (n_3759));
  AN22X1 g89901(.A (n_3170), .B (n_7022), .C (n_3171), .D (n_7020), .Q
       (n_3758));
  AN22X1 g89902(.A (n_3165), .B (n_6336), .C (n_3173), .D (n_6334), .Q
       (n_3757));
  AN22X1 g89903(.A (n_3170), .B (n_6340), .C (n_3171), .D (n_6338), .Q
       (n_3756));
  AO22X1 g89904(.A (n_3165), .B (n_7049), .C (n_3173), .D (n_7047), .Q
       (n_3755));
  AN22X1 g89906(.A (n_3171), .B (n_6307), .C (n_3165), .D (n_6305), .Q
       (n_3753));
  AN22X1 g89907(.A (n_3170), .B (n_6309), .C (n_3173), .D (n_6303), .Q
       (n_3752));
  NA2X1 g89909(.A (n_3341), .B (n_3340), .Q (n_3750));
  AN22X1 g89911(.A (n_3167), .B (n_7116), .C (n_2300), .D (n_7110), .Q
       (n_3748));
  AN22X1 g89912(.A (n_3167), .B (n_7023), .C (n_3177), .D (n_7021), .Q
       (n_3747));
  AN22X1 g89913(.A (n_3167), .B (n_6341), .C (n_3177), .D (n_6339), .Q
       (n_3746));
  AN22X1 g89914(.A (n_3167), .B (n_7054), .C (n_3177), .D (n_7052), .Q
       (n_3745));
  AN22X1 g89915(.A (n_3177), .B (n_6308), .C (n_3175), .D (n_6306), .Q
       (n_3744));
  AN22X1 g89916(.A (n_3167), .B (n_6310), .C (n_2300), .D (n_6304), .Q
       (n_3743));
  AN22X1 g89917(.A (n_3156), .B (n_6565), .C (n_3163), .D (n_6559), .Q
       (n_3742));
  AN22X1 g89918(.A (n_3152), .B (n_6902), .C (n_3163), .D (n_6900), .Q
       (n_3741));
  AN22X1 g89919(.A (n_3156), .B (n_6906), .C (n_3154), .D (n_6904), .Q
       (n_3740));
  AN22X1 g89920(.A (n_3152), .B (n_6406), .C (n_3163), .D (n_6404), .Q
       (n_3739));
  AN22X1 g89921(.A (n_3156), .B (n_6410), .C (n_3154), .D (n_6408), .Q
       (n_3738));
  AN22X1 g89922(.A (n_3154), .B (n_6563), .C (n_3152), .D (n_6561), .Q
       (n_3737));
  AN22X1 g89923(.A (n_3154), .B (n_6997), .C (n_3152), .D (n_6995), .Q
       (n_3736));
  AN22X1 g89924(.A (n_3156), .B (n_6999), .C (n_3163), .D (n_6993), .Q
       (n_3735));
  AN22X1 g89925(.A (n_3152), .B (n_6964), .C (n_3163), .D (n_6962), .Q
       (n_3734));
  AN22X1 g89926(.A (n_3156), .B (n_6968), .C (n_3154), .D (n_6966), .Q
       (n_3733));
  AN22X1 g89927(.A (n_3152), .B (n_6437), .C (n_3163), .D (n_6435), .Q
       (n_3732));
  AN22X1 g89928(.A (n_3156), .B (n_6441), .C (n_3154), .D (n_6439), .Q
       (n_3731));
  AN22X1 g89929(.A (n_3154), .B (n_6935), .C (n_3152), .D (n_6933), .Q
       (n_3730));
  AN22X1 g89930(.A (n_3156), .B (n_6937), .C (n_3163), .D (n_6931), .Q
       (n_3729));
  AN21X1 g89931(.A (n_3152), .B (n_7150), .C (n_3289), .Q (n_3728));
  AN21X1 g89932(.A (n_3156), .B (n_7154), .C (n_3288), .Q (n_3727));
  AN22X1 g89933(.A (n_3154), .B (n_7121), .C (n_3152), .D (n_7119), .Q
       (n_3726));
  AN22X1 g89934(.A (n_3156), .B (n_7123), .C (n_3163), .D (n_7117), .Q
       (n_3725));
  AN22X1 g89935(.A (n_3152), .B (n_7026), .C (n_3163), .D (n_7024), .Q
       (n_3724));
  AN22X1 g89936(.A (n_3156), .B (n_7030), .C (n_3154), .D (n_7028), .Q
       (n_3723));
  AN22X1 g89937(.A (n_3152), .B (n_6344), .C (n_3163), .D (n_6342), .Q
       (n_3722));
  AN22X1 g89938(.A (n_3156), .B (n_6348), .C (n_3154), .D (n_6346), .Q
       (n_3721));
  AN22X1 g89939(.A (n_3152), .B (n_7057), .C (n_3163), .D (n_7055), .Q
       (n_3720));
  AN22X1 g89940(.A (n_3156), .B (n_7061), .C (n_3154), .D (n_7059), .Q
       (n_3719));
  AN22X1 g89941(.A (n_3154), .B (n_6315), .C (n_3152), .D (n_6313), .Q
       (n_3718));
  AN22X1 g89942(.A (n_3156), .B (n_6317), .C (n_3163), .D (n_6311), .Q
       (n_3717));
  ON22X1 g89943(.A (n_3160), .B (n_2408), .C (n_3162), .D (n_2406), .Q
       (n_3716));
  ON22X1 g89944(.A (n_3160), .B (n_2410), .C (n_3162), .D (n_2446), .Q
       (n_3715));
  ON22X1 g89945(.A (n_3160), .B (n_2456), .C (n_3162), .D (n_2444), .Q
       (n_3714));
  AN22X1 g89946(.A (n_3159), .B (n_6965), .C (n_3161), .D (n_6963), .Q
       (n_3713));
  ON22X1 g89947(.A (n_3158), .B (n_2450), .C (n_3162), .D (n_2453), .Q
       (n_3712));
  AO22X1 g89948(.A (n_3159), .B (n_6934), .C (n_3161), .D (n_6932), .Q
       (n_3711));
  AN22X1 g89949(.A (n_3175), .B (n_7205), .C (n_2300), .D (n_7203), .Q
       (n_3710));
  AN221X1 g89950(.A (n_6667), .B (n_3073), .C (n_6672), .D (n_3052), .E
       (n_3129), .Q (n_3708));
  AN22X1 g89951(.A (n_3177), .B (n_6370), .C (n_3175), .D (n_6368), .Q
       (n_3707));
  NO2X1 g89952(.A (n_3308), .B (n_3309), .Q (n_3706));
  NO2X1 g89953(.A (n_3292), .B (n_3293), .Q (n_3705));
  AN22X1 g89954(.A (n_3167), .B (n_6372), .C (n_2300), .D (n_6366), .Q
       (n_3704));
  NO2X1 g89955(.A (n_3291), .B (n_3307), .Q (n_3703));
  NO2X1 g89956(.A (n_3290), .B (n_3383), .Q (n_3702));
  AN22X1 g89957(.A (n_3177), .B (n_7083), .C (n_3175), .D (n_7081), .Q
       (n_3701));
  AN22X1 g89958(.A (n_3167), .B (n_7085), .C (n_2300), .D (n_7079), .Q
       (n_3700));
  AN21X1 g89959(.A (n_3175), .B (n_6275), .C (n_3305), .Q (n_3699));
  AN22X1 g89960(.A (n_3167), .B (n_6279), .C (n_3177), .D (n_6277), .Q
       (n_3698));
  NA2X1 g89961(.A (n_3302), .B (n_3303), .Q (n_3697));
  NO2X1 g89963(.A (n_3300), .B (n_3301), .Q (n_3695));
  AN21X1 g89964(.A (n_3170), .B (n_7177), .C (n_3299), .Q (n_3694));
  NA2X1 g89965(.A (n_3297), .B (n_3298), .Q (n_3693));
  AO22X1 g89966(.A (n_3170), .B (n_6371), .C (n_3173), .D (n_6365), .Q
       (n_3692));
  NO2X1 g89967(.A (n_3295), .B (n_3296), .Q (n_3691));
  NO2X1 g89968(.A (n_3294), .B (n_3304), .Q (n_3690));
  AN22X1 g89969(.A (n_3171), .B (n_7082), .C (n_3165), .D (n_7080), .Q
       (n_3689));
  AN22X1 g89970(.A (n_3170), .B (n_7084), .C (n_3173), .D (n_7078), .Q
       (n_3688));
  AN22X1 g89971(.A (n_3165), .B (n_6274), .C (n_3173), .D (n_6272), .Q
       (n_3687));
  AN22X1 g89972(.A (n_3170), .B (n_6278), .C (n_3171), .D (n_6276), .Q
       (n_3686));
  AN221X1 g89973(.A (n_6357), .B (n_3073), .C (n_6358), .D (n_3075), .E
       (n_3228), .Q (n_3685));
  AN22X1 g89975(.A (n_3152), .B (n_7212), .C (n_3163), .D (n_7210), .Q
       (n_3683));
  AN22X1 g89976(.A (n_3156), .B (n_7216), .C (n_3154), .D (n_7214), .Q
       (n_3682));
  AN22X1 g89977(.A (n_3152), .B (n_6747), .C (n_3163), .D (n_6745), .Q
       (n_3681));
  AN22X1 g89978(.A (n_3156), .B (n_6751), .C (n_3154), .D (n_6749), .Q
       (n_3680));
  NA3X1 g89979(.A (n_3230), .B (n_3132), .C (n_3131), .Q (n_3679));
  AN22X1 g89980(.A (n_3154), .B (n_6377), .C (n_3152), .D (n_6375), .Q
       (n_3678));
  NO2X1 g89981(.A (n_3285), .B (n_3286), .Q (n_3677));
  AN21X1 g89982(.A (n_3156), .B (n_7185), .C (n_3284), .Q (n_3676));
  AN22X1 g89983(.A (n_3156), .B (n_6379), .C (n_3163), .D (n_6373), .Q
       (n_3675));
  NO2X1 g89987(.A (n_3282), .B (n_3283), .Q (n_3671));
  NO2X1 g89988(.A (n_3280), .B (n_3281), .Q (n_3670));
  AN221X1 g89989(.A (n_6326), .B (n_3073), .C (n_6327), .D (n_3075), .E
       (n_3145), .Q (n_3669));
  AN22X1 g89991(.A (n_3154), .B (n_7090), .C (n_3152), .D (n_7088), .Q
       (n_3667));
  AN22X1 g89992(.A (n_3156), .B (n_7092), .C (n_3163), .D (n_7086), .Q
       (n_3666));
  AN22X1 g89994(.A (n_3152), .B (n_6282), .C (n_3163), .D (n_6280), .Q
       (n_3664));
  AN22X1 g89995(.A (n_3156), .B (n_6286), .C (n_3154), .D (n_6284), .Q
       (n_3663));
  AN221X1 g89996(.A (n_7194), .B (n_3073), .C (n_7195), .D (n_3075), .E
       (n_3141), .Q (n_3662));
  NA2X1 g89997(.A (n_3264), .B (n_8561), .Q (n_3661));
  NA2X1 g89998(.A (n_3253), .B (n_3266), .Q (n_3660));
  AN22X1 g90000(.A (n_3157), .B (n_7122), .C (n_3159), .D (n_7120), .Q
       (n_3658));
  AO22X1 g90001(.A (n_3157), .B (n_6347), .C (n_3161), .D (n_6343), .Q
       (n_3657));
  AN22X1 g90003(.A (n_3159), .B (n_7151), .C (n_3161), .D (n_7149), .Q
       (n_3655));
  AN22X1 g90005(.A (n_3159), .B (n_7058), .C (n_3161), .D (n_7056), .Q
       (n_3653));
  NA2X1 g90006(.A (n_3242), .B (n_3252), .Q (n_3652));
  NO2X2 g90007(.A (n_3250), .B (n_3239), .Q (n_3651));
  ON21X1 g90010(.A (n_3162), .B (n_2461), .C (n_2640), .Q (n_3648));
  AN22X1 g90011(.A (n_3175), .B (n_6709), .C (n_2300), .D (n_6707), .Q
       (n_3647));
  AN22X1 g90012(.A (n_3167), .B (n_6713), .C (n_3177), .D (n_6711), .Q
       (n_3646));
  AN22X1 g90015(.A (n_3165), .B (n_6708), .C (n_3173), .D (n_6706), .Q
       (n_3643));
  AN22X1 g90016(.A (n_3170), .B (n_6712), .C (n_3171), .D (n_6710), .Q
       (n_3642));
  AN22X1 g90017(.A (n_3165), .B (n_6677), .C (n_3173), .D (n_6675), .Q
       (n_3641));
  AN22X1 g90018(.A (n_3170), .B (n_6681), .C (n_3171), .D (n_6679), .Q
       (n_3640));
  AN22X1 g90019(.A (n_3157), .B (n_6750), .C (n_3161), .D (n_6746), .Q
       (n_3639));
  AO22X1 g90020(.A (n_3157), .B (n_6378), .C (n_3159), .D (n_6376), .Q
       (n_3638));
  AN22X1 g90022(.A (n_3157), .B (n_6285), .C (n_3161), .D (n_6281), .Q
       (n_3636));
  ON22X1 g90023(.A (n_3158), .B (n_2451), .C (n_2586), .D (n_2407), .Q
       (n_3635));
  ON22X1 g90024(.A (n_3158), .B (n_2449), .C (n_2586), .D (n_2452), .Q
       (n_3634));
  ON22X1 g90025(.A (n_3158), .B (n_2448), .C (n_2586), .D (n_2411), .Q
       (n_3633));
  AN22X1 g90026(.A (n_3157), .B (n_6967), .C (n_2587), .D (n_6969), .Q
       (n_3632));
  ON22X1 g90027(.A (n_3158), .B (n_2402), .C (n_2586), .D (n_2403), .Q
       (n_3631));
  NO2X1 g90029(.A (n_3272), .B (n_3273), .Q (n_3629));
  AN22X1 g90030(.A (n_3159), .B (n_7089), .C (n_3161), .D (n_7087), .Q
       (n_3628));
  ON22X1 g90032(.A (n_3160), .B (n_2454), .C (n_2586), .D (n_2409), .Q
       (n_3626));
  AN22X1 g90033(.A (n_3175), .B (n_6802), .C (n_2300), .D (n_6800), .Q
       (n_3625));
  AN22X1 g90034(.A (n_3167), .B (n_6806), .C (n_3177), .D (n_6804), .Q
       (n_3624));
  AO22X1 g90035(.A (n_3175), .B (n_6833), .C (n_2300), .D (n_6831), .Q
       (n_3623));
  AO22X1 g90036(.A (n_3167), .B (n_6837), .C (n_3177), .D (n_6835), .Q
       (n_3622));
  AN22X1 g90037(.A (n_3175), .B (n_6771), .C (n_2300), .D (n_6769), .Q
       (n_3621));
  AN22X1 g90038(.A (n_3167), .B (n_6775), .C (n_3177), .D (n_6773), .Q
       (n_3620));
  AN22X1 g90041(.A (n_3175), .B (n_6864), .C (n_2300), .D (n_6862), .Q
       (n_3617));
  AN22X1 g90042(.A (n_3167), .B (n_6868), .C (n_3177), .D (n_6866), .Q
       (n_3616));
  AN22X1 g90043(.A (n_3167), .B (n_7209), .C (n_3177), .D (n_7207), .Q
       (n_3615));
  AN22X1 g90044(.A (n_3165), .B (n_6801), .C (n_3173), .D (n_6799), .Q
       (n_3614));
  AN22X1 g90045(.A (n_3170), .B (n_6805), .C (n_3171), .D (n_6803), .Q
       (n_3613));
  AN22X1 g90046(.A (n_3165), .B (n_6832), .C (n_3173), .D (n_6830), .Q
       (n_3612));
  AN22X1 g90047(.A (n_3170), .B (n_6836), .C (n_3171), .D (n_6834), .Q
       (n_3611));
  AN22X1 g90048(.A (n_3165), .B (n_6770), .C (n_3173), .D (n_6768), .Q
       (n_3610));
  AN22X1 g90049(.A (n_3170), .B (n_6774), .C (n_3171), .D (n_6772), .Q
       (n_3609));
  AN22X1 g90050(.A (n_3170), .B (n_6526), .C (n_3171), .D (n_6524), .Q
       (n_3608));
  NO2X1 g90051(.A (n_3243), .B (n_3245), .Q (n_3607));
  AN22X1 g90052(.A (n_3165), .B (n_6863), .C (n_3173), .D (n_6861), .Q
       (n_3606));
  AN22X1 g90053(.A (n_3170), .B (n_6867), .C (n_3171), .D (n_6865), .Q
       (n_3605));
  AN22X1 g90054(.A (n_3152), .B (n_6716), .C (n_3163), .D (n_6714), .Q
       (n_3604));
  AN22X1 g90055(.A (n_3156), .B (n_6720), .C (n_3154), .D (n_6718), .Q
       (n_3603));
  AN22X1 g90056(.A (n_3152), .B (n_6685), .C (n_3163), .D (n_6683), .Q
       (n_3602));
  AN22X1 g90057(.A (n_3156), .B (n_6689), .C (n_3154), .D (n_6687), .Q
       (n_3601));
  AN221X1 g90058(.A (n_6691), .B (n_3066), .C (n_6703), .D (n_3052), .E
       (n_3130), .Q (n_3600));
  AN22X1 g90059(.A (n_3152), .B (n_6809), .C (n_3163), .D (n_6807), .Q
       (n_3599));
  AN22X1 g90060(.A (n_3156), .B (n_6813), .C (n_3154), .D (n_6811), .Q
       (n_3598));
  AN22X1 g90061(.A (n_3152), .B (n_6840), .C (n_3163), .D (n_6838), .Q
       (n_3597));
  AN22X1 g90062(.A (n_3156), .B (n_6844), .C (n_3154), .D (n_6842), .Q
       (n_3596));
  AN22X1 g90063(.A (n_3154), .B (n_6780), .C (n_3152), .D (n_6778), .Q
       (n_3595));
  AN22X1 g90064(.A (n_3156), .B (n_6782), .C (n_3163), .D (n_6776), .Q
       (n_3594));
  AN22X1 g90065(.A (n_3152), .B (n_6530), .C (n_3163), .D (n_6528), .Q
       (n_3593));
  AN22X1 g90067(.A (n_3152), .B (n_6871), .C (n_3163), .D (n_6869), .Q
       (n_3591));
  AN22X1 g90068(.A (n_3156), .B (n_6875), .C (n_3154), .D (n_6873), .Q
       (n_3590));
  AN221X1 g90069(.A (n_6791), .B (n_3073), .C (n_6796), .D (n_3052), .E
       (n_3127), .Q (n_3589));
  AN222X1 g90070(.A (n_3073), .B (n_6822), .C (n_6823), .D (n_3075), .E
       (n_6827), .F (n_3051), .Q (n_3588));
  AN221X1 g90071(.A (n_6760), .B (n_3073), .C (n_6765), .D (n_3052), .E
       (n_3126), .Q (n_3587));
  AN22X1 g90074(.A (n_3157), .B (n_7153), .C (n_2587), .D (n_7155), .Q
       (n_3584));
  AO22X2 g90075(.A (n_3157), .B (n_7029), .C (n_2587), .D (n_7031), .Q
       (n_3583));
  AN22X1 g90076(.A (n_3157), .B (n_7060), .C (n_2587), .D (n_7062), .Q
       (n_3582));
  AN22X1 g90077(.A (n_3161), .B (n_7118), .C (n_2587), .D (n_7124), .Q
       (n_3581));
  ON22X1 g90078(.A (n_3162), .B (n_2404), .C (n_2586), .D (n_2405), .Q
       (n_3580));
  AO22X2 g90079(.A (n_3159), .B (n_6345), .C (n_2587), .D (n_6349), .Q
       (n_3579));
  AN221X1 g90080(.A (n_6605), .B (n_3073), .C (n_6599), .D (n_3107), .E
       (n_3113), .Q (n_3578));
  ON22X1 g90082(.A (n_3158), .B (n_2455), .C (n_2586), .D (n_2445), .Q
       (n_3576));
  AN22X1 g90084(.A (n_3157), .B (n_7091), .C (n_2587), .D (n_7093), .Q
       (n_3574));
  AO22X2 g90085(.A (n_3161), .B (n_6374), .C (n_2587), .D (n_6380), .Q
       (n_3573));
  AN22X1 g90086(.A (n_3159), .B (n_6748), .C (n_2587), .D (n_6752), .Q
       (n_3572));
  AN22X1 g90088(.A (n_3159), .B (n_6283), .C (n_2587), .D (n_6287), .Q
       (n_3570));
  AN22X1 g90091(.A (n_3157), .B (n_6719), .C (n_3161), .D (n_6715), .Q
       (n_3567));
  AN22X1 g90092(.A (n_3157), .B (n_6688), .C (n_3161), .D (n_6684), .Q
       (n_3566));
  AN22X1 g90093(.A (n_3157), .B (n_6812), .C (n_3161), .D (n_6808), .Q
       (n_3565));
  AN22X1 g90094(.A (n_3159), .B (n_6841), .C (n_3161), .D (n_6839), .Q
       (n_3564));
  AO22X2 g90095(.A (n_3159), .B (n_6779), .C (n_3161), .D (n_6777), .Q
       (n_3563));
  AO22X2 g90096(.A (n_3157), .B (n_6533), .C (n_3161), .D (n_6529), .Q
       (n_3562));
  AN22X1 g90097(.A (n_3157), .B (n_6874), .C (n_3161), .D (n_6870), .Q
       (n_3561));
  AO22X1 g90098(.A (n_3167), .B (n_6620), .C (n_3177), .D (n_6618), .Q
       (n_3560));
  AN22X1 g90099(.A (n_3171), .B (n_6493), .C (n_3177), .D (n_6494), .Q
       (n_3559));
  AO22X1 g90100(.A (n_3170), .B (n_6495), .C (n_3167), .D (n_6496), .Q
       (n_3558));
  AO22X1 g90101(.A (n_3167), .B (n_6465), .C (n_3177), .D (n_6463), .Q
       (n_3557));
  AN22X1 g90102(.A (n_3159), .B (n_6717), .C (n_2587), .D (n_6721), .Q
       (n_3556));
  AN22X1 g90103(.A (n_3159), .B (n_6686), .C (n_2587), .D (n_6690), .Q
       (n_3555));
  AO22X1 g90104(.A (n_3165), .B (n_6460), .C (n_3173), .D (n_6458), .Q
       (n_3554));
  AO22X1 g90105(.A (n_3175), .B (n_6616), .C (n_2300), .D (n_6614), .Q
       (n_3553));
  AN22X1 g90106(.A (n_3165), .B (n_6615), .C (n_3173), .D (n_6613), .Q
       (n_3552));
  AN22X1 g90107(.A (n_3170), .B (n_6619), .C (n_3171), .D (n_6617), .Q
       (n_3551));
  AO22X2 g90108(.A (n_3177), .B (n_6587), .C (n_3175), .D (n_6585), .Q
       (n_3550));
  AO22X1 g90109(.A (n_3167), .B (n_6589), .C (n_2300), .D (n_6583), .Q
       (n_3549));
  AN22X1 g90110(.A (n_3171), .B (n_6586), .C (n_3165), .D (n_6584), .Q
       (n_3548));
  AN22X1 g90111(.A (n_3170), .B (n_6588), .C (n_3173), .D (n_6582), .Q
       (n_3547));
  AN22X1 g90112(.A (n_3165), .B (n_6491), .C (n_3175), .D (n_6492), .Q
       (n_3546));
  AO22X2 g90113(.A (n_3173), .B (n_6489), .C (n_2300), .D (n_6490), .Q
       (n_3545));
  AO22X1 g90114(.A (n_3175), .B (n_6461), .C (n_2300), .D (n_6459), .Q
       (n_3544));
  AO22X1 g90115(.A (n_3170), .B (n_6464), .C (n_3171), .D (n_6462), .Q
       (n_3543));
  AN22X1 g90116(.A (n_3159), .B (n_6810), .C (n_2587), .D (n_6814), .Q
       (n_3542));
  AN22X1 g90117(.A (n_3157), .B (n_6843), .C (n_2587), .D (n_6845), .Q
       (n_3541));
  AO22X1 g90118(.A (n_3157), .B (n_6781), .C (n_2587), .D (n_6783), .Q
       (n_3540));
  NA2X2 g90119(.A (n_3235), .B (n_2611), .Q (n_3539));
  AN22X1 g90120(.A (n_3159), .B (n_6872), .C (n_2587), .D (n_6876), .Q
       (n_3538));
  AN22X1 g90121(.A (n_3152), .B (n_6592), .C (n_3163), .D (n_6590), .Q
       (n_3537));
  AN22X1 g90122(.A (n_3152), .B (n_6499), .C (n_3163), .D (n_6497), .Q
       (n_3536));
  AN22X1 g90123(.A (n_3152), .B (n_6468), .C (n_3163), .D (n_6466), .Q
       (n_3535));
  AN22X1 g90124(.A (n_3156), .B (n_6596), .C (n_3154), .D (n_6594), .Q
       (n_3534));
  AN22X1 g90125(.A (n_3156), .B (n_6503), .C (n_3154), .D (n_6501), .Q
       (n_3533));
  AN22X1 g90126(.A (n_3156), .B (n_6472), .C (n_3154), .D (n_6470), .Q
       (n_3532));
  AN22X1 g90127(.A (n_3156), .B (n_6627), .C (n_2340), .D (n_6608), .Q
       (n_3531));
  AO22X1 g90128(.A (n_3154), .B (n_6625), .C (n_3157), .D (n_6626), .Q
       (n_3530));
  AN22X1 g90129(.A (n_3163), .B (n_6621), .C (n_3161), .D (n_6622), .Q
       (n_3529));
  AN22X1 g90130(.A (n_3152), .B (n_6623), .C (n_3159), .D (n_6624), .Q
       (n_3528));
  AN22X1 g90131(.A (n_3157), .B (n_6595), .C (n_3161), .D (n_6591), .Q
       (n_3527));
  AN22X1 g90132(.A (n_3157), .B (n_6502), .C (n_3161), .D (n_6498), .Q
       (n_3526));
  ON22X1 g90133(.A (n_3160), .B (n_2397), .C (n_3162), .D (n_2394), .Q
       (n_3525));
  AN22X1 g90134(.A (n_3159), .B (n_6500), .C (n_2587), .D (n_6504), .Q
       (n_3524));
  AN22X1 g90135(.A (n_3159), .B (n_6593), .C (n_2587), .D (n_6597), .Q
       (n_3523));
  NO2X1 g90136(.A (n_3007), .B (n_3179), .Q (n_3709));
  INX1 g90138(.A (n_2346), .Q (csr_data_out[25]));
  NA2X1 g90139(.A (n_2678), .B (csr_data_out[15]), .Q (n_3522));
  ON21X1 g90140(.A (n_2533), .B (n_2590), .C (csr_data_out[14]), .Q
       (n_3521));
  ON21X1 g90142(.A (n_2535), .B (n_2590), .C (csr_data_out[13]), .Q
       (n_3520));
  ON21X1 g90143(.A (n_2527), .B (n_2590), .C (csr_data_out[12]), .Q
       (n_3519));
  ON21X1 g90144(.A (n_2529), .B (n_2590), .C (csr_data_out[6]), .Q
       (n_3518));
  OA21X2 g90145(.A (n_2526), .B (n_2590), .C (csr_data_out[8]), .Q
       (n_3517));
  NO2I1X4 g90146(.B (n_2715), .AN (csr_data_out[2]), .Q (n_3516));
  OA21X4 g90147(.A (n_2576), .B (n_2646), .C (csr_data_out[4]), .Q
       (n_3515));
  ON21X1 g90148(.A (n_2524), .B (n_2590), .C (csr_data_out[9]), .Q
       (n_3514));
  NA2X2 g90149(.A (n_2651), .B (csr_data_out[5]), .Q (n_3513));
  AN22X1 g90150(.A (n_3104), .B (n_6359), .C (n_3055), .D (n_6356), .Q
       (n_3512));
  AN22X1 g90151(.A (n_3104), .B (n_6731), .C (n_3055), .D (n_6728), .Q
       (n_3511));
  AO22X1 g90152(.A (n_3104), .B (n_7196), .C (n_3055), .D (n_7193), .Q
       (n_3510));
  AN22X1 g90153(.A (n_3054), .B (n_7200), .C (n_3063), .D (n_7201), .Q
       (n_3509));
  AN22X1 g90154(.A (n_3105), .B (n_6268), .C (n_2339), .D (n_6267), .Q
       (n_3508));
  AN22X1 g90155(.A (n_3054), .B (n_6270), .C (n_3063), .D (n_6271), .Q
       (n_3507));
  AN22X1 g90156(.A (n_3105), .B (n_7074), .C (n_2339), .D (n_7073), .Q
       (n_3506));
  AN22X1 g90157(.A (n_3054), .B (n_7076), .C (n_3063), .D (n_7077), .Q
       (n_3505));
  AN22X1 g90158(.A (n_3063), .B (n_6643), .C (n_3105), .D (n_6640), .Q
       (n_3504));
  AN22X1 g90159(.A (n_3105), .B (n_7167), .C (n_2339), .D (n_7166), .Q
       (n_3503));
  AN22X1 g90160(.A (n_3054), .B (n_7169), .C (n_3063), .D (n_7170), .Q
       (n_3502));
  AO22X1 g90161(.A (n_3105), .B (n_6361), .C (n_2339), .D (n_6360), .Q
       (n_3501));
  AN22X1 g90162(.A (n_3054), .B (n_6363), .C (n_3063), .D (n_6364), .Q
       (n_3500));
  AN22X1 g90163(.A (n_3105), .B (n_6733), .C (n_2340), .D (n_6732), .Q
       (n_3499));
  AN22X1 g90164(.A (n_3054), .B (n_6735), .C (n_3063), .D (n_6736), .Q
       (n_3498));
  AN22X1 g90166(.A (n_3054), .B (n_6921), .C (n_3051), .D (n_6920), .Q
       (n_3496));
  NO2X1 g90167(.A (n_3213), .B (n_3215), .Q (n_3495));
  AN22X1 g90168(.A (n_3061), .B (n_6384), .C (n_2336), .D (n_6383), .Q
       (n_3494));
  AN21X1 g90169(.A (n_2336), .B (n_6538), .C (n_3209), .Q (n_3493));
  AN21X1 g90170(.A (n_3059), .B (n_6972), .C (n_3206), .Q (n_3492));
  NA2X1 g90171(.A (n_3193), .B (n_3205), .Q (n_3491));
  NO2X1 g90172(.A (n_3204), .B (n_3192), .Q (n_3490));
  AN21X1 g90173(.A (n_2336), .B (n_6879), .C (n_3201), .Q (n_3489));
  ON22X1 g90174(.A (n_3062), .B (n_2400), .C (n_2335), .D (n_2401), .Q
       (n_3488));
  AN22X1 g90175(.A (n_3057), .B (n_6386), .C (n_3064), .D (n_6385), .Q
       (n_3487));
  AN21X1 g90176(.A (n_3057), .B (n_6541), .C (n_3208), .Q (n_3486));
  AN22X1 g90177(.A (n_3057), .B (n_6975), .C (n_3064), .D (n_6974), .Q
       (n_3485));
  AO22X1 g90178(.A (n_3057), .B (n_6417), .C (n_3064), .D (n_6416), .Q
       (n_3484));
  NO2X1 g90179(.A (n_3202), .B (n_3231), .Q (n_3483));
  AN21X1 g90180(.A (n_3057), .B (n_6882), .C (n_3199), .Q (n_3482));
  AN21X1 g90182(.A (n_2336), .B (n_7220), .C (n_3214), .Q (n_3480));
  AN21X1 g90183(.A (n_3104), .B (n_7227), .C (n_3212), .Q (n_3479));
  AN21X1 g90184(.A (n_2339), .B (n_7228), .C (n_3198), .Q (n_3478));
  AN22X1 g90185(.A (n_3054), .B (n_7231), .C (n_3063), .D (n_7232), .Q
       (n_3477));
  AN22X1 g90186(.A (n_3104), .B (n_6545), .C (n_3055), .D (n_6542), .Q
       (n_3476));
  AN22X1 g90187(.A (n_3104), .B (n_6421), .C (n_3055), .D (n_6418), .Q
       (n_3475));
  AN21X1 g90188(.A (n_3104), .B (n_6886), .C (n_3200), .Q (n_3474));
  AN22X1 g90189(.A (n_3104), .B (n_6390), .C (n_3055), .D (n_6387), .Q
       (n_3473));
  AN21X1 g90190(.A (n_3104), .B (n_6979), .C (n_3195), .Q (n_3472));
  AN21X1 g90191(.A (n_3104), .B (n_6948), .C (n_3194), .Q (n_3471));
  AN22X1 g90192(.A (n_3104), .B (n_6917), .C (n_3055), .D (n_6914), .Q
       (n_3470));
  AN22X1 g90193(.A (n_3107), .B (n_7219), .C (n_3069), .D (n_7218), .Q
       (n_3469));
  AN22X1 g90194(.A (n_3105), .B (n_6888), .C (n_2340), .D (n_6887), .Q
       (n_3468));
  AN22X1 g90196(.A (n_3105), .B (n_6392), .C (n_2339), .D (n_6391), .Q
       (n_3466));
  AN22X1 g90197(.A (n_3054), .B (n_6549), .C (n_3063), .D (n_6550), .Q
       (n_3465));
  AN21X1 g90198(.A (n_2339), .B (n_6546), .C (n_3188), .Q (n_3464));
  AN22X1 g90199(.A (n_3063), .B (n_6984), .C (n_3073), .D (n_6977), .Q
       (n_3463));
  AN22X1 g90200(.A (n_3054), .B (n_6425), .C (n_3063), .D (n_6426), .Q
       (n_3462));
  AN22X1 g90201(.A (n_3105), .B (n_6981), .C (n_2339), .D (n_6980), .Q
       (n_3461));
  AN22X1 g90202(.A (n_3054), .B (n_6952), .C (n_3063), .D (n_6953), .Q
       (n_3460));
  AN22X1 g90203(.A (n_3105), .B (n_6423), .C (n_2340), .D (n_6422), .Q
       (n_3459));
  AN21X1 g90204(.A (n_2339), .B (n_6949), .C (n_3187), .Q (n_3458));
  AN22X1 g90205(.A (n_3054), .B (n_6890), .C (n_3063), .D (n_6891), .Q
       (n_3457));
  AN22X1 g90206(.A (n_3063), .B (n_6922), .C (n_3073), .D (n_6915), .Q
       (n_3456));
  AN22X1 g90207(.A (n_3105), .B (n_6919), .C (n_2339), .D (n_6918), .Q
       (n_3455));
  AN22X1 g90208(.A (n_3057), .B (n_7130), .C (n_3064), .D (n_7129), .Q
       (n_3454));
  AN22X1 g90209(.A (n_3057), .B (n_7099), .C (n_3064), .D (n_7098), .Q
       (n_3453));
  AN22X1 g90210(.A (n_3057), .B (n_7006), .C (n_3064), .D (n_7005), .Q
       (n_3452));
  AN22X1 g90211(.A (n_3057), .B (n_6324), .C (n_3064), .D (n_6323), .Q
       (n_3451));
  AN22X1 g90212(.A (n_3057), .B (n_7037), .C (n_3064), .D (n_7036), .Q
       (n_3450));
  AO22X1 g90213(.A (n_3057), .B (n_6293), .C (n_3064), .D (n_6292), .Q
       (n_3449));
  AO22X1 g90217(.A (n_3073), .B (n_6946), .C (n_3075), .D (n_6947), .Q
       (n_3445));
  AN22X1 g90218(.A (n_3057), .B (n_7192), .C (n_3064), .D (n_7191), .Q
       (n_3444));
  AN22X1 g90220(.A (n_3057), .B (n_6355), .C (n_3064), .D (n_6354), .Q
       (n_3442));
  AO22X1 g90221(.A (n_3057), .B (n_7161), .C (n_3064), .D (n_7160), .Q
       (n_3441));
  AN22X1 g90222(.A (n_3057), .B (n_7068), .C (n_3064), .D (n_7067), .Q
       (n_3440));
  AN22X1 g90223(.A (n_3057), .B (n_6634), .C (n_3064), .D (n_6633), .Q
       (n_3439));
  AN22X1 g90224(.A (n_3057), .B (n_6262), .C (n_3064), .D (n_6261), .Q
       (n_3438));
  AO22X1 g90225(.A (n_3107), .B (n_6382), .C (n_2337), .D (n_6381), .Q
       (n_3437));
  AN22X1 g90226(.A (n_3107), .B (n_6537), .C (n_3069), .D (n_6536), .Q
       (n_3436));
  AN22X1 g90227(.A (n_3107), .B (n_6413), .C (n_3069), .D (n_6412), .Q
       (n_3435));
  AN22X1 g90228(.A (n_3107), .B (n_6940), .C (n_3071), .D (n_6939), .Q
       (n_3434));
  AN22X1 g90229(.A (n_3107), .B (n_6878), .C (n_3069), .D (n_6877), .Q
       (n_3433));
  AN21X1 g90230(.A (n_3059), .B (n_7127), .C (n_3186), .Q (n_3432));
  AN22X1 g90231(.A (n_3104), .B (n_7134), .C (n_3055), .D (n_7131), .Q
       (n_3431));
  AN22X1 g90233(.A (n_3104), .B (n_7103), .C (n_3055), .D (n_7100), .Q
       (n_3429));
  AN22X1 g90234(.A (n_3061), .B (n_7004), .C (n_2336), .D (n_7003), .Q
       (n_3428));
  AN22X1 g90235(.A (n_3104), .B (n_7010), .C (n_3055), .D (n_7007), .Q
       (n_3427));
  AN22X1 g90236(.A (n_3061), .B (n_6322), .C (n_3059), .D (n_6321), .Q
       (n_3426));
  AN22X1 g90238(.A (n_3061), .B (n_7035), .C (n_3059), .D (n_7034), .Q
       (n_3424));
  AN22X1 g90239(.A (n_3104), .B (n_7041), .C (n_2339), .D (n_7042), .Q
       (n_3423));
  AO22X2 g90240(.A (n_3061), .B (n_6291), .C (n_2336), .D (n_6290), .Q
       (n_3422));
  AN22X1 g90241(.A (n_3104), .B (n_6297), .C (n_3055), .D (n_6294), .Q
       (n_3421));
  AN22X1 g90242(.A (n_3054), .B (n_7138), .C (n_3063), .D (n_7139), .Q
       (n_3420));
  AN22X1 g90243(.A (n_3105), .B (n_7136), .C (n_2339), .D (n_7135), .Q
       (n_3419));
  AN22X1 g90244(.A (n_3054), .B (n_7107), .C (n_3063), .D (n_7108), .Q
       (n_3418));
  NA2X1 g90245(.A (n_3227), .B (n_3224), .Q (n_3417));
  AN22X1 g90246(.A (n_3054), .B (n_7014), .C (n_3063), .D (n_7015), .Q
       (n_3416));
  AN22X1 g90247(.A (n_3105), .B (n_7012), .C (n_2339), .D (n_7011), .Q
       (n_3415));
  AN22X1 g90248(.A (n_3054), .B (n_6332), .C (n_3063), .D (n_6333), .Q
       (n_3414));
  NA2X1 g90249(.A (n_3226), .B (n_3225), .Q (n_3413));
  AN22X1 g90250(.A (n_3063), .B (n_7046), .C (n_3105), .D (n_7043), .Q
       (n_3412));
  AN22X1 g90251(.A (n_3054), .B (n_6301), .C (n_3063), .D (n_6302), .Q
       (n_3411));
  AN22X1 g90252(.A (n_3105), .B (n_6299), .C (n_2339), .D (n_6298), .Q
       (n_3410));
  AN22X1 g90253(.A (n_3054), .B (n_6983), .C (n_3051), .D (n_6982), .Q
       (n_3409));
  AO22X1 g90255(.A (n_3061), .B (n_6725), .C (n_3059), .D (n_6724), .Q
       (n_3407));
  AO22X2 g90256(.A (n_3061), .B (n_6353), .C (n_3059), .D (n_6352), .Q
       (n_3406));
  AN22X1 g90257(.A (n_3061), .B (n_7066), .C (n_3059), .D (n_7065), .Q
       (n_3405));
  AO22X1 g90258(.A (n_3061), .B (n_7159), .C (n_3060), .D (n_7158), .Q
       (n_3404));
  AN22X1 g90259(.A (n_3061), .B (n_6632), .C (n_2336), .D (n_6631), .Q
       (n_3403));
  AN22X1 g90260(.A (n_3061), .B (n_6260), .C (n_3059), .D (n_6259), .Q
       (n_3402));
  AN22X1 g90261(.A (n_3061), .B (n_7190), .C (n_2336), .D (n_7189), .Q
       (n_3401));
  AN21X1 g90262(.A (n_3107), .B (n_7126), .C (n_3140), .Q (n_3400));
  AN22X1 g90263(.A (n_3107), .B (n_7095), .C (n_2337), .D (n_7094), .Q
       (n_3399));
  AN22X1 g90264(.A (n_3107), .B (n_7002), .C (n_2337), .D (n_7001), .Q
       (n_3398));
  AN22X1 g90265(.A (n_3107), .B (n_6320), .C (n_3071), .D (n_6319), .Q
       (n_3397));
  AN22X1 g90266(.A (n_3107), .B (n_7033), .C (n_2337), .D (n_7032), .Q
       (n_3396));
  AN22X1 g90267(.A (n_3107), .B (n_6289), .C (n_3071), .D (n_6288), .Q
       (n_3395));
  NO2I1X1 g90269(.B (n_3151), .AN (n_6924), .Q (n_3393));
  NO2I1X1 g90270(.B (n_3176), .AN (n_6926), .Q (n_3392));
  NO2I1X1 g90271(.B (n_3151), .AN (n_6986), .Q (n_3391));
  NO2I1X1 g90272(.B (n_3178), .AN (n_6990), .Q (n_3390));
  NO2I1X1 g90273(.B (n_3176), .AN (n_6988), .Q (n_3389));
  NO2I1X1 g90274(.B (n_3151), .AN (n_6955), .Q (n_3388));
  NO2I1X1 g90275(.B (n_3174), .AN (n_6923), .Q (n_3387));
  NO2I1X1 g90276(.B (n_3174), .AN (n_6985), .Q (n_3386));
  NO2I1X1 g90277(.B (n_3166), .AN (n_6987), .Q (n_3385));
  NA3X1 g90278(.A (n_2957), .B (n_3096), .C (n_3015), .Q
       (csr_data_out[11]));
  NA3X1 g90279(.A (n_2950), .B (n_3023), .C (n_3089), .Q
       (csr_data_out[16]));
  NA3X1 g90280(.A (n_3211), .B (n_2884), .C (n_2862), .Q
       (csr_data_out[17]));
  NA3X1 g90281(.A (n_3217), .B (n_2863), .C (n_2848), .Q
       (csr_data_out[18]));
  NA3X1 g90282(.A (n_2949), .B (n_3025), .C (n_3090), .Q
       (csr_data_out[20]));
  NA3X1 g90283(.A (n_3216), .B (n_2865), .C (n_2873), .Q
       (csr_data_out[23]));
  NA3X1 g90284(.A (n_2967), .B (n_3028), .C (n_3091), .Q
       (csr_data_out[19]));
  NA3X1 g90285(.A (n_2954), .B (n_3027), .C (n_3092), .Q
       (csr_data_out[21]));
  NA3X1 g90286(.A (n_2956), .B (n_3029), .C (n_3093), .Q
       (csr_data_out[24]));
  NA3X1 g90287(.A (n_3099), .B (n_3088), .C (n_2928), .Q
       (csr_data_out[7]));
  NA3X1 g90289(.A (n_3221), .B (n_2885), .C (n_2874), .Q
       (csr_data_out[27]));
  NA3X1 g90290(.A (n_3220), .B (n_2875), .C (n_2879), .Q
       (csr_data_out[28]));
  NA3X1 g90291(.A (n_3222), .B (n_2876), .C (n_2877), .Q
       (csr_data_out[29]));
  NA3X1 g90292(.A (n_2958), .B (n_3095), .C (n_3030), .Q
       (csr_data_out[31]));
  NA3X1 g90293(.A (n_2959), .B (n_3097), .C (n_3034), .Q
       (csr_data_out[26]));
  NA3X1 g90294(.A (n_3223), .B (n_2882), .C (n_2880), .Q
       (csr_data_out[30]));
  NA3X1 g90295(.A (n_2960), .B (n_3098), .C (n_3036), .Q
       (csr_data_out[22]));
  NO2I1X1 g90296(.B (n_3151), .AN (n_6645), .Q (n_3383));
  AN22X1 g90297(.A (n_3104), .B (n_6638), .C (n_3055), .D (n_6635), .Q
       (n_3382));
  AN22X1 g90298(.A (n_3104), .B (n_6266), .C (n_3055), .D (n_6263), .Q
       (n_3381));
  AN22X1 g90299(.A (n_3104), .B (n_7072), .C (n_3055), .D (n_7069), .Q
       (n_3380));
  AN21X1 g90300(.A (n_3107), .B (n_6723), .C (n_3138), .Q (n_3379));
  AN22X1 g90301(.A (n_3107), .B (n_6351), .C (n_2337), .D (n_6350), .Q
       (n_3378));
  NO2X1 g90303(.A (n_3147), .B (n_3135), .Q (n_3376));
  AN21X1 g90304(.A (n_3107), .B (n_7064), .C (n_3137), .Q (n_3375));
  AN22X1 g90305(.A (n_3107), .B (n_6258), .C (n_2337), .D (n_6257), .Q
       (n_3374));
  AN22X1 g90306(.A (n_3107), .B (n_7188), .C (n_3071), .D (n_7187), .Q
       (n_3373));
  AN22X1 g90312(.A (n_3057), .B (n_6696), .C (n_3064), .D (n_6695), .Q
       (n_3367));
  AN22X1 g90313(.A (n_3104), .B (n_6700), .C (n_3055), .D (n_6697), .Q
       (n_3366));
  AN22X1 g90314(.A (n_3057), .B (n_6665), .C (n_3064), .D (n_6664), .Q
       (n_3365));
  AN22X1 g90315(.A (n_3104), .B (n_6669), .C (n_3055), .D (n_6666), .Q
       (n_3364));
  AN22X1 g90316(.A (n_3054), .B (n_7045), .C (n_3051), .D (n_7044), .Q
       (n_3363));
  AN22X1 g90317(.A (n_3054), .B (n_6704), .C (n_3107), .D (n_6692), .Q
       (n_3362));
  AN22X1 g90318(.A (n_3052), .B (n_6641), .C (n_3107), .D (n_6630), .Q
       (n_3361));
  AN22X1 g90320(.A (n_3061), .B (n_6694), .C (n_3059), .D (n_6693), .Q
       (n_3360));
  AN22X1 g90321(.A (n_3061), .B (n_6663), .C (n_3059), .D (n_6662), .Q
       (n_3359));
  AN22X1 g90322(.A (n_3105), .B (n_6702), .C (n_2339), .D (n_6701), .Q
       (n_3358));
  AN22X1 g90323(.A (n_3105), .B (n_6671), .C (n_2339), .D (n_6670), .Q
       (n_3357));
  AN22X1 g90324(.A (n_3107), .B (n_6785), .C (n_3064), .D (n_6788), .Q
       (n_3356));
  AN22X1 g90325(.A (n_3104), .B (n_6793), .C (n_3055), .D (n_6790), .Q
       (n_3355));
  AN22X1 g90326(.A (n_3057), .B (n_6820), .C (n_3064), .D (n_6819), .Q
       (n_3354));
  AN22X1 g90327(.A (n_3104), .B (n_6824), .C (n_3055), .D (n_6821), .Q
       (n_3353));
  AN22X1 g90328(.A (n_3057), .B (n_6758), .C (n_3064), .D (n_6757), .Q
       (n_3352));
  AN22X1 g90329(.A (n_3104), .B (n_6762), .C (n_3055), .D (n_6759), .Q
       (n_3351));
  AN22X1 g90330(.A (n_3057), .B (n_6510), .C (n_3064), .D (n_6509), .Q
       (n_3350));
  AN22X1 g90331(.A (n_3104), .B (n_6514), .C (n_3055), .D (n_6511), .Q
       (n_3349));
  AN22X1 g90332(.A (n_3057), .B (n_6851), .C (n_3064), .D (n_6850), .Q
       (n_3348));
  AN22X1 g90333(.A (n_3104), .B (n_6855), .C (n_3055), .D (n_6852), .Q
       (n_3347));
  AN22X1 g90334(.A (n_3054), .B (n_6673), .C (n_3063), .D (n_6674), .Q
       (n_3346));
  NO2I1X1 g90335(.B (n_3160), .AN (n_7244), .Q (n_3345));
  NO2I1X1 g90336(.B (n_3158), .AN (n_7246), .Q (n_3344));
  NA2X1 g90339(.A (n_3177), .B (n_7145), .Q (n_3341));
  NA2X1 g90340(.A (n_3167), .B (n_7147), .Q (n_3340));
  NA2X1 g90343(.A (n_3173), .B (n_6737), .Q (n_3338));
  NA2X1 g90344(.A (n_3165), .B (n_6739), .Q (n_3337));
  NA2X1 g90345(.A (n_3173), .B (n_7140), .Q (n_3336));
  NA2X1 g90346(.A (n_3165), .B (n_7142), .Q (n_3335));
  AO22X1 g90350(.A (n_3073), .B (n_6264), .C (n_3075), .D (n_6265), .Q
       (n_3331));
  AN22X1 g90351(.A (n_3061), .B (n_6787), .C (n_3060), .D (n_6786), .Q
       (n_3330));
  AN22X1 g90352(.A (n_3061), .B (n_6818), .C (n_3059), .D (n_6817), .Q
       (n_3329));
  AN22X1 g90353(.A (n_3061), .B (n_6756), .C (n_2336), .D (n_6755), .Q
       (n_3328));
  AN22X1 g90354(.A (n_3061), .B (n_6508), .C (n_3060), .D (n_6507), .Q
       (n_3327));
  AN22X1 g90355(.A (n_3061), .B (n_6849), .C (n_3060), .D (n_6848), .Q
       (n_3326));
  AN22X1 g90356(.A (n_3105), .B (n_6795), .C (n_2339), .D (n_6794), .Q
       (n_3325));
  AN22X1 g90357(.A (n_3105), .B (n_6826), .C (n_2339), .D (n_6825), .Q
       (n_3324));
  AN22X1 g90358(.A (n_3105), .B (n_6764), .C (n_2340), .D (n_6763), .Q
       (n_3323));
  AN22X1 g90359(.A (n_3105), .B (n_6516), .C (n_2339), .D (n_6515), .Q
       (n_3322));
  AN22X1 g90360(.A (n_3105), .B (n_6857), .C (n_2339), .D (n_6856), .Q
       (n_3321));
  AN22X1 g90361(.A (n_3054), .B (n_6797), .C (n_3063), .D (n_6798), .Q
       (n_3320));
  AN22X1 g90363(.A (n_3054), .B (n_6766), .C (n_3063), .D (n_6767), .Q
       (n_3318));
  AN22X1 g90364(.A (n_3054), .B (n_6518), .C (n_3063), .D (n_6519), .Q
       (n_3317));
  AN22X1 g90365(.A (n_3054), .B (n_6859), .C (n_3063), .D (n_6860), .Q
       (n_3316));
  AN22X1 g90366(.A (n_3107), .B (n_6661), .C (n_2337), .D (n_6660), .Q
       (n_3315));
  NO2I1X1 g90367(.B (n_3162), .AN (n_6994), .Q (n_3314));
  NA2X1 g90368(.A (n_3159), .B (n_6996), .Q (n_3313));
  NA2X1 g90369(.A (n_3157), .B (n_6998), .Q (n_3312));
  AN22X1 g90370(.A (n_3057), .B (n_6789), .C (n_2337), .D (n_6784), .Q
       (n_3311));
  AN22X1 g90371(.A (n_3107), .B (n_6754), .C (n_2337), .D (n_6753), .Q
       (n_3310));
  NO2I1X1 g90372(.B (n_3151), .AN (n_7172), .Q (n_3309));
  NO2I1X1 g90373(.B (n_3176), .AN (n_7174), .Q (n_3308));
  NO2I1X1 g90374(.B (n_3176), .AN (n_6647), .Q (n_3307));
  AN22X1 g90375(.A (n_3104), .B (n_7165), .C (n_3055), .D (n_7162), .Q
       (n_3306));
  NO2I1X1 g90376(.B (n_3151), .AN (n_6273), .Q (n_3305));
  NO2I1X1 g90377(.B (n_3174), .AN (n_6644), .Q (n_3304));
  NA2X1 g90378(.A (n_3173), .B (n_7202), .Q (n_3303));
  NA2X1 g90379(.A (n_3165), .B (n_7204), .Q (n_3302));
  NO2I1X1 g90380(.B (n_3174), .AN (n_7171), .Q (n_3301));
  NO2I1X1 g90381(.B (n_3166), .AN (n_7173), .Q (n_3300));
  NO2I1X1 g90382(.B (n_3172), .AN (n_7175), .Q (n_3299));
  NA2X1 g90383(.A (n_3165), .B (n_6367), .Q (n_3298));
  NA2X1 g90384(.A (n_3171), .B (n_6369), .Q (n_3297));
  NO2I1X1 g90385(.B (n_3166), .AN (n_6646), .Q (n_3296));
  NO2I1X1 g90386(.B (n_3172), .AN (n_6648), .Q (n_3295));
  NO2I1X1 g90387(.B (n_3169), .AN (n_6650), .Q (n_3294));
  NO2I1X1 g90388(.B (n_3178), .AN (n_7176), .Q (n_3293));
  NO2I1X1 g90389(.B (n_3168), .AN (n_7178), .Q (n_3292));
  NO2I1X1 g90390(.B (n_3178), .AN (n_6649), .Q (n_3291));
  NO2I1X1 g90391(.B (n_3168), .AN (n_6651), .Q (n_3290));
  NO2I1X1 g90392(.B (n_3164), .AN (n_7148), .Q (n_3289));
  NO2I1X1 g90393(.B (n_3155), .AN (n_7152), .Q (n_3288));
  AN22X1 g90394(.A (n_3063), .B (n_6705), .C (n_3073), .D (n_6698), .Q
       (n_3287));
  NO2I1X1 g90395(.B (n_3164), .AN (n_7179), .Q (n_3286));
  NO2I1X1 g90396(.B (n_3153), .AN (n_7181), .Q (n_3285));
  NO2I1X1 g90397(.B (n_3155), .AN (n_7183), .Q (n_3284));
  NO2I1X1 g90398(.B (n_3153), .AN (n_6654), .Q (n_3283));
  NO2I1X1 g90399(.B (n_3155), .AN (n_6656), .Q (n_3282));
  NO2I1X1 g90400(.B (n_3164), .AN (n_6652), .Q (n_3281));
  NO2I1X1 g90401(.B (n_2280), .AN (n_6658), .Q (n_3280));
  AO22X2 g90404(.A (n_3107), .B (n_6816), .C (n_3071), .D (n_6815), .Q
       (n_3277));
  AN22X1 g90405(.A (n_3107), .B (n_6506), .C (n_2337), .D (n_6505), .Q
       (n_3276));
  AN22X1 g90406(.A (n_3107), .B (n_6847), .C (n_2337), .D (n_6846), .Q
       (n_3275));
  NO2I1X1 g90408(.B (n_3158), .AN (n_7184), .Q (n_3274));
  NO2I1X1 g90409(.B (n_3162), .AN (n_6653), .Q (n_3273));
  NO2I1X1 g90410(.B (n_3160), .AN (n_6655), .Q (n_3272));
  AN22X1 g90411(.A (n_3063), .B (n_6612), .C (n_3105), .D (n_6609), .Q
       (n_3271));
  AN22X1 g90412(.A (n_3054), .B (n_6580), .C (n_3063), .D (n_6581), .Q
       (n_3270));
  AN22X1 g90414(.A (n_3054), .B (n_6456), .C (n_3063), .D (n_6457), .Q
       (n_3268));
  AO22X1 g90415(.A (n_3061), .B (n_6601), .C (n_3060), .D (n_6600), .Q
       (n_3267));
  AN22X1 g90416(.A (n_3057), .B (n_6603), .C (n_3064), .D (n_6602), .Q
       (n_3266));
  AN22X1 g90418(.A (n_3057), .B (n_6572), .C (n_3064), .D (n_6571), .Q
       (n_3264));
  AN22X1 g90419(.A (n_3057), .B (n_6479), .C (n_3064), .D (n_6478), .Q
       (n_3263));
  AN22X1 g90420(.A (n_3061), .B (n_6446), .C (n_3059), .D (n_6445), .Q
       (n_3262));
  AN22X1 g90421(.A (n_3057), .B (n_6448), .C (n_3064), .D (n_6447), .Q
       (n_3261));
  AN22X1 g90422(.A (n_3061), .B (n_6477), .C (n_3060), .D (n_6476), .Q
       (n_3260));
  NO2I1X1 g90423(.B (n_3151), .AN (n_6676), .Q (n_3259));
  NO2I1X1 g90425(.B (n_3178), .AN (n_6680), .Q (n_3257));
  AN22X1 g90427(.A (n_3107), .B (n_6568), .C (n_3069), .D (n_6567), .Q
       (n_3255));
  NA2X1 g90428(.A (n_3115), .B (n_3119), .Q (n_3254));
  AN22X1 g90429(.A (n_3104), .B (n_6607), .C (n_3055), .D (n_6604), .Q
       (n_3253));
  AN22X1 g90430(.A (n_3104), .B (n_6576), .C (n_3055), .D (n_6573), .Q
       (n_3252));
  ON22X1 g90431(.A (n_3103), .B (n_2392), .C (n_3056), .D (n_2393), .Q
       (n_3251));
  AO22X1 g90432(.A (n_3104), .B (n_6452), .C (n_3055), .D (n_6449), .Q
       (n_3250));
  AND2X1 g90434(.A (n_3167), .B (n_6527), .Q (n_3248));
  AND2X2 g90436(.A (n_3177), .B (n_6525), .Q (n_3247));
  NO2I1X1 g90437(.B (n_3176), .AN (n_6523), .Q (n_3246));
  NO2I1X1 g90438(.B (n_3174), .AN (n_6520), .Q (n_3245));
  NO2I1X1 g90440(.B (n_3166), .AN (n_6522), .Q (n_3243));
  AN22X1 g90441(.A (n_3105), .B (n_6578), .C (n_2340), .D (n_6577), .Q
       (n_3242));
  NA2X1 g90442(.A (n_3123), .B (n_3112), .Q (n_3241));
  AN22X1 g90443(.A (n_3107), .B (n_6444), .C (n_2337), .D (n_6443), .Q
       (n_3240));
  NA2X1 g90444(.A (n_3150), .B (n_3114), .Q (n_3239));
  ON22X1 g90445(.A (n_3074), .B (n_2398), .C (n_3076), .D (n_2399), .Q
       (n_3238));
  ON22X1 g90446(.A (n_3074), .B (n_2395), .C (n_3076), .D (n_2396), .Q
       (n_3237));
  AO22X2 g90447(.A (n_3073), .B (n_6481), .C (n_3075), .D (n_6482), .Q
       (n_3236));
  NA2X1 g90448(.A (n_3159), .B (n_6531), .Q (n_3235));
  AN22X1 g90449(.A (n_3054), .B (n_6611), .C (n_3052), .D (n_6610), .Q
       (n_3234));
  AN22X1 g90450(.A (n_3066), .B (n_6598), .C (n_2587), .D (n_6628), .Q
       (n_3233));
  NO2I1X1 g90451(.B (n_3158), .AN (n_6471), .Q (n_3232));
  NA2X1 g90452(.A (n_3182), .B (n_7275), .Q (n_3384));
  NA3X1 g90453(.A (n_2999), .B (n_3101), .C (n_2979), .Q
       (csr_data_out[3]));
  NO2I1X1 g90454(.B (n_3065), .AN (n_6943), .Q (n_3231));
  NO2X1 g90455(.A (n_8563), .B (n_2758), .Q (n_7860));
  NO2X1 g90456(.A (n_8563), .B (n_2596), .Q (n_7859));
  NA2X1 g90457(.A (n_3051), .B (n_7168), .Q (n_3230));
  NO2X1 g90459(.A (n_2281), .B (n_2447), .Q (n_3228));
  NA2X1 g90460(.A (n_3105), .B (n_7105), .Q (n_3227));
  NA2X1 g90461(.A (n_3105), .B (n_6330), .Q (n_3226));
  NA2X1 g90462(.A (n_2339), .B (n_6329), .Q (n_3225));
  NA2X1 g90463(.A (n_2339), .B (n_7104), .Q (n_3224));
  AN211X1 g90464(.A (n_2731), .B (csr_mtvec[30]), .C (n_3010), .D
       (n_3035), .Q (n_3223));
  AN211X1 g90465(.A (n_2731), .B (csr_mtvec[29]), .C (n_3039), .D
       (n_3031), .Q (n_3222));
  AN211X1 g90466(.A (n_2731), .B (csr_mtvec[27]), .C (n_3002), .D
       (n_3032), .Q (n_3221));
  AN211X1 g90467(.A (n_2731), .B (csr_mtvec[28]), .C (n_3041), .D
       (n_3033), .Q (n_3220));
  NO2I1X1 g90469(.B (n_2338), .AN (n_6908), .Q (n_3218));
  AND4X1 g90470(.A (n_2987), .B (n_2830), .C (n_2932), .D (n_2773), .Q
       (n_3217));
  AND4X1 g90471(.A (n_2832), .B (n_2929), .C (n_2990), .D (n_2774), .Q
       (n_3216));
  NO2I1X1 g90472(.B (n_3065), .AN (n_7222), .Q (n_3215));
  NO2I1X1 g90473(.B (n_3062), .AN (n_7221), .Q (n_3214));
  NO2I1X1 g90474(.B (n_3058), .AN (n_7223), .Q (n_3213));
  NO2I1X1 g90475(.B (n_3056), .AN (n_7224), .Q (n_3212));
  AN211X1 g90476(.A (n_2731), .B (csr_mtvec[17]), .C (n_2983), .D
       (n_3024), .Q (n_3211));
  NO2I1X1 g90477(.B (n_2281), .AN (n_6889), .Q (n_3210));
  NO2I1X1 g90478(.B (n_3062), .AN (n_6539), .Q (n_3209));
  NO2I1X1 g90479(.B (n_3065), .AN (n_6540), .Q (n_3208));
  NO2I1X1 g90481(.B (n_3062), .AN (n_6973), .Q (n_3206));
  NA2X1 g90482(.A (n_3061), .B (n_6415), .Q (n_3205));
  NO2I1X1 g90483(.B (n_3062), .AN (n_6942), .Q (n_3204));
  OR2X1 g90484(.A (n_3109), .B (n_2316), .Q (n_3203));
  NO2I1X1 g90485(.B (n_3058), .AN (n_6944), .Q (n_3202));
  NO2I1X1 g90486(.B (n_3062), .AN (n_6880), .Q (n_3201));
  NO2I1X1 g90487(.B (n_3056), .AN (n_6883), .Q (n_3200));
  NO2I1X1 g90488(.B (n_3065), .AN (n_6881), .Q (n_3199));
  NO2I1X1 g90489(.B (n_3106), .AN (n_7229), .Q (n_3198));
  NO2I1X1 g90491(.B (n_2281), .AN (n_7230), .Q (n_3196));
  NO2I1X1 g90492(.B (n_3056), .AN (n_6976), .Q (n_3195));
  NO2I1X1 g90493(.B (n_3056), .AN (n_6945), .Q (n_3194));
  NA2X1 g90494(.A (n_2336), .B (n_6414), .Q (n_3193));
  NO2I1X1 g90495(.B (n_2335), .AN (n_6941), .Q (n_3192));
  NO2I1X1 g90496(.B (n_3108), .AN (n_6971), .Q (n_3191));
  NO2I1X1 g90497(.B (n_3108), .AN (n_6909), .Q (n_3190));
  NO2I1X1 g90499(.B (n_3106), .AN (n_6547), .Q (n_3188));
  NO2I1X1 g90500(.B (n_3106), .AN (n_6950), .Q (n_3187));
  NO2I1X1 g90501(.B (n_3062), .AN (n_7128), .Q (n_3186));
  NA3X1 g90503(.A (n_2948), .B (n_3016), .C (n_3000), .Q
       (csr_data_out[10]));
  NA3X1 g90504(.A (n_3100), .B (n_2823), .C (n_2972), .Q
       (csr_data_out[4]));
  NA3X2 g90505(.A (n_3017), .B (n_2980), .C (n_2978), .Q
       (csr_data_out[2]));
  NA3X1 g90506(.A (n_2962), .B (n_2997), .C (n_2981), .Q
       (csr_data_out[6]));
  NA3X1 g90507(.A (n_3094), .B (n_2985), .C (n_2841), .Q
       (csr_data_out[8]));
  NA3X1 g90508(.A (n_2955), .B (n_3011), .C (n_2995), .Q
       (csr_data_out[9]));
  NA3X1 g90509(.A (n_2963), .B (n_2977), .C (n_2973), .Q
       (csr_data_out[5]));
  NA3X1 g90510(.A (n_2951), .B (n_3021), .C (n_3014), .Q
       (csr_data_out[15]));
  NA3X1 g90511(.A (n_2952), .B (n_3020), .C (n_3013), .Q
       (csr_data_out[13]));
  NA3X1 g90512(.A (n_3037), .B (n_3022), .C (n_3012), .Q
       (csr_data_out[12]));
  NA3X1 g90513(.A (n_2953), .B (n_3026), .C (n_3018), .Q
       (csr_data_out[14]));
  NO2X1 g90514(.A (n_8563), .B (n_2815), .Q (n_8297));
  INX6 g90516(.A (n_3178), .Q (n_3177));
  INX8 g90517(.A (n_3176), .Q (n_3175));
  INX6 g90518(.A (n_3174), .Q (n_3173));
  INX4 g90519(.A (n_3172), .Q (n_3171));
  INX8 g90520(.A (n_3169), .Q (n_3170));
  INX6 g90521(.A (n_3168), .Q (n_3167));
  INX8 g90522(.A (n_3166), .Q (n_3165));
  INX4 g90523(.A (n_3164), .Q (n_3163));
  INX6 g90524(.A (n_3162), .Q (n_3161));
  INX8 g90525(.A (n_3160), .Q (n_3159));
  INX8 g90526(.A (n_3158), .Q (n_3157));
  INX6 g90527(.A (n_2280), .Q (n_3156));
  INX8 g90528(.A (n_3155), .Q (n_3154));
  INX6 g90529(.A (n_3153), .Q (n_3152));
  NA2X1 g90531(.A (n_3105), .B (n_6454), .Q (n_3150));
  NO2I1X1 g90532(.B (n_2281), .AN (n_6393), .Q (n_3149));
  NO2I1X1 g90534(.B (n_3053), .AN (n_6642), .Q (n_3147));
  NO2I1X1 g90536(.B (n_2281), .AN (n_6331), .Q (n_3145));
  NO2I1X1 g90539(.B (n_2281), .AN (n_6951), .Q (n_3142));
  NO2I1X1 g90540(.B (n_2281), .AN (n_7199), .Q (n_3141));
  NO2I1X1 g90541(.B (n_2338), .AN (n_7125), .Q (n_3140));
  NO2I1X1 g90543(.B (n_2338), .AN (n_6722), .Q (n_3138));
  NO2I1X1 g90544(.B (n_2338), .AN (n_7063), .Q (n_3137));
  NO2I1X1 g90546(.B (n_2338), .AN (n_6629), .Q (n_3135));
  AND2X1 g90547(.A (n_3052), .B (n_6517), .Q (n_3134));
  NO2I1X1 g90548(.B (n_2281), .AN (n_6858), .Q (n_3133));
  NA2X1 g90549(.A (n_3075), .B (n_7164), .Q (n_3132));
  NA2X1 g90550(.A (n_3073), .B (n_7163), .Q (n_3131));
  NO2I1X1 g90551(.B (n_3076), .AN (n_6699), .Q (n_3130));
  NO2I1X1 g90552(.B (n_3076), .AN (n_6668), .Q (n_3129));
  NO2I1X1 g90554(.B (n_3076), .AN (n_6792), .Q (n_3127));
  NO2I1X1 g90555(.B (n_3076), .AN (n_6761), .Q (n_3126));
  NA2X1 g90558(.A (n_3105), .B (n_6485), .Q (n_3123));
  NA2X1 g90562(.A (n_3107), .B (n_6475), .Q (n_3119));
  NO2I1X1 g90564(.B (n_3062), .AN (n_6570), .Q (n_3118));
  AND2X1 g90565(.A (n_3052), .B (n_6486), .Q (n_3117));
  NA2X1 g90567(.A (n_2340), .B (n_6484), .Q (n_3115));
  NA2X1 g90568(.A (n_2340), .B (n_6453), .Q (n_3114));
  NO2I1X1 g90569(.B (n_3076), .AN (n_6606), .Q (n_3113));
  NA2X1 g90570(.A (n_3066), .B (n_6474), .Q (n_3112));
  OR2X1 g90571(.A (n_3077), .B (n_2504), .Q (n_3184));
  OR2X1 g90572(.A (n_3077), .B (n_2602), .Q (n_3183));
  NA2X1 g90573(.A (n_3050), .B (n_2944), .Q (n_3182));
  OR2X1 g90574(.A (n_3078), .B (n_2504), .Q (n_3181));
  OR2X1 g90575(.A (n_3078), .B (n_2602), .Q (n_3180));
  OA21X1 g90576(.A (n_3045), .B (n_2442), .C (n_8300), .Q (n_3179));
  OR2X4 g90577(.A (n_3081), .B (n_2851), .Q (n_3178));
  OR2X4 g90578(.A (n_3081), .B (n_2856), .Q (n_3176));
  OR2X4 g90579(.A (n_3080), .B (n_2853), .Q (n_3174));
  OR2X4 g90580(.A (n_3080), .B (n_2851), .Q (n_3172));
  OR2X4 g90581(.A (n_3080), .B (n_2857), .Q (n_3169));
  OR2X4 g90582(.A (n_3081), .B (n_2857), .Q (n_3168));
  OR2X4 g90583(.A (n_3080), .B (n_2856), .Q (n_3166));
  NA2X4 g90584(.A (n_3082), .B (n_2854), .Q (n_3164));
  OR3X4 g90585(.A (n_3005), .B (n_2917), .C (n_2853), .Q (n_3162));
  NA2X4 g90586(.A (n_3049), .B (n_2328), .Q (n_3160));
  OR3X4 g90587(.A (n_2917), .B (n_3005), .C (n_2851), .Q (n_3158));
  NA2X4 g90589(.A (n_3082), .B (n_2850), .Q (n_3155));
  NA2X4 g90590(.A (n_3082), .B (n_2328), .Q (n_3153));
  OR2X4 g90591(.A (n_3081), .B (n_2853), .Q (n_3151));
  BUX8 g90595(.A (n_2340), .Q (n_2339));
  INX8 g90597(.A (n_3108), .Q (n_3107));
  INX8 g90598(.A (n_3106), .Q (n_3105));
  INX8 g90599(.A (n_3103), .Q (n_3104));
  OR2X1 g90601(.A (n_3043), .B (n_3042), .Q (n_3102));
  AN221X1 g90602(.A (csr_mcause[3]), .B (n_2725), .C (n_7964), .D
       (n_2323), .E (n_8565), .Q (n_3101));
  AN221X1 g90603(.A (csr_mscratch[4]), .B (n_2727), .C (n_7892), .D
       (n_2323), .E (n_2986), .Q (n_3100));
  AN221X1 g90604(.A (csr_mcause[7]), .B (n_2725), .C (n_7923), .D
       (n_2323), .E (n_2992), .Q (n_3099));
  AN21X1 g90605(.A (n_2731), .B (csr_mtvec[22]), .C (n_3019), .Q
       (n_3098));
  AN21X1 g90606(.A (n_2731), .B (csr_mtvec[26]), .C (n_3009), .Q
       (n_3097));
  AN211X1 g90607(.A (n_2324), .B (n_4433), .C (n_2822), .D (n_2993), .Q
       (n_3096));
  AN21X1 g90608(.A (n_2731), .B (csr_mtvec[31]), .C (n_3038), .Q
       (n_3095));
  AN221X1 g90609(.A (csr_mscratch[8]), .B (n_2727), .C (n_7895), .D
       (n_2323), .E (n_3001), .Q (n_3094));
  AN21X1 g90610(.A (n_2731), .B (csr_mtvec[24]), .C (n_2991), .Q
       (n_3093));
  AN21X1 g90611(.A (n_2731), .B (csr_mtvec[21]), .C (n_2996), .Q
       (n_3092));
  AN21X1 g90612(.A (n_2731), .B (csr_mtvec[19]), .C (n_2989), .Q
       (n_3091));
  AN21X1 g90613(.A (n_2731), .B (csr_mtvec[20]), .C (n_2988), .Q
       (n_3090));
  AN21X1 g90614(.A (n_2731), .B (csr_mtvec[16]), .C (n_2982), .Q
       (n_3089));
  AN221X1 g90615(.A (n_4434), .B (n_2324), .C (n_8029), .D (n_2735), .E
       (n_2994), .Q (n_3088));
  ON21X1 g90616(.A (n_2945), .B (n_7714), .C (n_2503), .Q (n_8206));
  AO21X1 g90618(.A (n_8165), .B (n_2626), .C (n_3042), .Q (n_3110));
  ON21X1 g90619(.A (n_7708), .B (n_2627), .C (n_2969), .Q (n_3109));
  NO2X4 g90620(.A (n_2937), .B (n_3005), .Q (n_2340));
  NA2X4 g90621(.A (n_2938), .B (n_2334), .Q (n_3108));
  NA2X4 g90622(.A (n_2939), .B (n_2332), .Q (n_3106));
  NA2X4 g90623(.A (n_2938), .B (n_2332), .Q (n_3103));
  INX8 g90624(.A (n_3076), .Q (n_3075));
  INX8 g90625(.A (n_3074), .Q (n_3073));
  INX2 g90627(.A (n_2338), .Q (n_3071));
  INX2 g90629(.A (n_2338), .Q (n_3069));
  INX4 g90632(.A (n_2338), .Q (n_2337));
  INX8 g90635(.A (n_3066), .Q (n_2338));
  INX6 g90636(.A (n_3065), .Q (n_3064));
  INX8 g90637(.A (n_3048), .Q (n_3063));
  INX8 g90638(.A (n_3062), .Q (n_3061));
  BUX2 g90639(.A (n_3060), .Q (n_3059));
  INX3 g90643(.A (n_2335), .Q (n_2336));
  INX6 g90645(.A (n_3058), .Q (n_3057));
  INX6 g90646(.A (n_3056), .Q (n_3055));
  INX6 g90647(.A (n_3053), .Q (n_3054));
  BUX6 g90649(.A (n_3052), .Q (n_3051));
  AND6X1 g90651(.A (n_2946), .B (n_2704), .C (n_2705), .D (n_2925), .E
       (n_2706), .F (n_2702), .Q (n_3050));
  NA2X1 g90652(.A (n_3047), .B (n_2504), .Q (n_3087));
  NA2X1 g90653(.A (n_3046), .B (n_2504), .Q (n_3086));
  NA2X1 g90654(.A (n_3046), .B (n_2602), .Q (n_3085));
  NA2X1 g90655(.A (n_3047), .B (n_2602), .Q (n_3084));
  AND2X2 g90656(.A (n_2333), .B (n_2330), .Q (n_3049));
  NA2X1 g90657(.A (n_3047), .B (n_2805), .Q (n_3083));
  NA2X1 g90658(.A (n_3045), .B (n_2442), .Q (n_8300));
  AND2X4 g90659(.A (n_2332), .B (n_2330), .Q (n_3082));
  NA2X4 g90660(.A (n_3004), .B (n_2330), .Q (n_3081));
  NA2X4 g90661(.A (n_2334), .B (n_2330), .Q (n_3080));
  NA2X1 g90662(.A (n_3046), .B (n_2805), .Q (n_3079));
  NA2X1 g90663(.A (n_3046), .B (n_2804), .Q (n_3078));
  NA2X1 g90664(.A (n_3047), .B (n_2804), .Q (n_3077));
  NA2X4 g90665(.A (n_2942), .B (n_2333), .Q (n_3076));
  NA2X4 g90666(.A (n_2942), .B (n_2332), .Q (n_3074));
  NO2X4 g90667(.A (n_2943), .B (n_3003), .Q (n_3066));
  NA2X4 g90668(.A (n_2939), .B (n_3004), .Q (n_3065));
  NA2X2 g90669(.A (n_2936), .B (n_2333), .Q (n_3048));
  NA2X4 g90670(.A (n_2939), .B (n_2334), .Q (n_3062));
  NO2X4 g90671(.A (n_2937), .B (n_3003), .Q (n_3060));
  NA2X4 g90672(.A (n_2936), .B (n_2334), .Q (n_3058));
  NA2X4 g90673(.A (n_2936), .B (n_3004), .Q (n_3056));
  NA2X4 g90674(.A (n_2936), .B (n_2332), .Q (n_3053));
  NO2X4 g90675(.A (n_2940), .B (n_3005), .Q (n_3052));
  INX1 g90677(.A (n_3047), .Q (n_3046));
  HAX1 g90678(.A (n_2802), .B (n_2440), .S (n_3047), .CO (n_3045));
  AO222X1 g90679(.A (n_8046), .B (n_2735), .C (csr_mcycle[28]), .D
       (n_2755), .E (csr_minstret[28]), .F (n_2733), .Q (n_3041));
  NO2X1 g90680(.A (n_8165), .B (n_2481), .Q (n_3040));
  AO222X1 g90681(.A (n_8047), .B (n_2735), .C (csr_mcycle[29]), .D
       (n_2755), .E (csr_minstret[29]), .F (n_2733), .Q (n_3039));
  AO222X1 g90682(.A (n_8049), .B (n_2735), .C (csr_mcycle[63]), .D
       (n_2756), .E (csr_minstret[63]), .F (n_2732), .Q (n_3038));
  AN211X1 g90683(.A (n_2727), .B (csr_mscratch[12]), .C (n_2849), .D
       (n_2871), .Q (n_3037));
  AN221X1 g90684(.A (csr_mcycle[54]), .B (n_2756), .C
       (csr_minstret[54]), .D (n_2732), .E (n_2843), .Q (n_3036));
  ON211X1 g90685(.A (n_2325), .B (n_4450), .C (n_2934), .D (n_2825), .Q
       (n_3035));
  AN221X1 g90686(.A (csr_mcycle[58]), .B (n_2756), .C
       (csr_minstret[58]), .D (n_2732), .E (n_2840), .Q (n_3034));
  NA2X1 g90687(.A (n_2922), .B (n_2839), .Q (n_3033));
  NA2X1 g90688(.A (n_2966), .B (n_2836), .Q (n_3032));
  NA2X1 g90689(.A (n_2965), .B (n_2837), .Q (n_3031));
  AN221X1 g90690(.A (csr_mcycle[31]), .B (n_2755), .C
       (csr_minstret[31]), .D (n_2733), .E (n_2838), .Q (n_3030));
  AN221X1 g90691(.A (csr_mcycle[56]), .B (n_2756), .C
       (csr_minstret[56]), .D (n_2732), .E (n_2829), .Q (n_3029));
  AN221X1 g90692(.A (csr_mcycle[51]), .B (n_2756), .C
       (csr_minstret[51]), .D (n_2732), .E (n_2828), .Q (n_3028));
  AN221X1 g90693(.A (csr_mcycle[53]), .B (n_2756), .C
       (csr_minstret[53]), .D (n_2732), .E (n_2833), .Q (n_3027));
  AN222X1 g90694(.A (n_2756), .B (csr_mcycle[46]), .C
       (csr_minstret[46]), .D (n_2732), .E (n_7902), .F (n_2323), .Q
       (n_3026));
  AN221X1 g90695(.A (csr_mcycle[52]), .B (n_2756), .C
       (csr_minstret[52]), .D (n_2732), .E (n_2831), .Q (n_3025));
  NA2X1 g90696(.A (n_2930), .B (n_2827), .Q (n_3024));
  AN221X1 g90697(.A (csr_mcycle[48]), .B (n_2756), .C
       (csr_minstret[48]), .D (n_2732), .E (n_2826), .Q (n_3023));
  AN222X1 g90698(.A (n_2756), .B (csr_mcycle[44]), .C
       (csr_minstret[44]), .D (n_2732), .E (csr_mtval[12]), .F
       (n_2726), .Q (n_3022));
  AN222X1 g90699(.A (n_2756), .B (csr_mcycle[47]), .C
       (csr_minstret[47]), .D (n_2732), .E (csr_mtval[15]), .F
       (n_2726), .Q (n_3021));
  AN222X1 g90700(.A (n_2756), .B (csr_mcycle[45]), .C
       (csr_minstret[45]), .D (n_2732), .E (csr_mtval[13]), .F
       (n_2726), .Q (n_3020));
  AO222X1 g90701(.A (n_8039), .B (n_2735), .C (csr_mcycle[22]), .D
       (n_2755), .E (csr_minstret[22]), .F (n_2733), .Q (n_3019));
  AN222X1 g90702(.A (n_2755), .B (csr_mcycle[14]), .C
       (csr_minstret[14]), .D (n_2733), .E (csr_mtvec[14]), .F
       (n_2731), .Q (n_3018));
  AN221X1 g90703(.A (csr_mcause[2]), .B (n_2725), .C (n_7890), .D
       (n_2323), .E (n_2931), .Q (n_3017));
  AN222X1 g90704(.A (n_2756), .B (csr_mcycle[42]), .C
       (csr_minstret[42]), .D (n_2732), .E (n_7897), .F (n_2323), .Q
       (n_3016));
  AN222X1 g90705(.A (n_2756), .B (csr_mcycle[43]), .C
       (csr_minstret[43]), .D (n_2732), .E (csr_mtvec[11]), .F
       (n_2731), .Q (n_3015));
  AN222X1 g90706(.A (n_2755), .B (csr_mcycle[15]), .C
       (csr_minstret[15]), .D (n_2733), .E (csr_mtvec[15]), .F
       (n_2731), .Q (n_3014));
  AN222X1 g90707(.A (n_2755), .B (csr_mcycle[13]), .C
       (csr_minstret[13]), .D (n_2733), .E (csr_mtvec[13]), .F
       (n_2731), .Q (n_3013));
  AN222X1 g90708(.A (n_2755), .B (csr_mcycle[12]), .C
       (csr_minstret[12]), .D (n_2733), .E (csr_mtvec[12]), .F
       (n_2731), .Q (n_3012));
  AN222X0 g90709(.A (n_2756), .B (csr_mcycle[41]), .C
       (csr_minstret[41]), .D (n_2732), .E (n_7896), .F (n_2323), .Q
       (n_3011));
  AO222X1 g90710(.A (n_8048), .B (n_2735), .C (csr_mcycle[30]), .D
       (n_2755), .E (csr_minstret[30]), .F (n_2733), .Q (n_3010));
  AO222X1 g90711(.A (n_8043), .B (n_2735), .C (csr_mcycle[26]), .D
       (n_2755), .E (csr_minstret[26]), .F (n_2733), .Q (n_3009));
  AND2X1 g90712(.A (n_2945), .B (n_2571), .Q (n_3008));
  OR2X1 g90713(.A (n_7707), .B (n_2627), .Q (n_3044));
  NO2X1 g90714(.A (n_7710), .B (n_2627), .Q (n_3043));
  AO21X1 g90715(.A (n_957), .B (n_2635), .C (n_2316), .Q (n_3042));
  INX1 g90716(.A (n_3006), .Q (n_3007));
  INX4 g90721(.A (n_2333), .Q (n_3005));
  INX2 g90724(.A (n_3004), .Q (n_3003));
  AO222X1 g90727(.A (n_8045), .B (n_2735), .C (csr_mcycle[27]), .D
       (n_2755), .E (csr_minstret[27]), .F (n_2733), .Q (n_3002));
  NA2X1 g90728(.A (n_2927), .B (n_2819), .Q (n_3001));
  AN222X1 g90729(.A (n_2755), .B (csr_mcycle[10]), .C
       (csr_minstret[10]), .D (n_2733), .E (csr_mtvec[10]), .F
       (n_2731), .Q (n_3000));
  AN211X1 g90730(.A (n_2727), .B (csr_mscratch[3]), .C (n_2818), .D
       (n_2820), .Q (n_2999));
  AN222X1 g90731(.A (n_2755), .B (csr_mcycle[25]), .C
       (csr_minstret[25]), .D (n_2733), .E (n_8042), .F (n_2735), .Q
       (n_2998));
  AN222X1 g90732(.A (n_2756), .B (csr_mcycle[38]), .C
       (csr_minstret[38]), .D (n_2732), .E (n_7894), .F (n_2323), .Q
       (n_2997));
  AO222X1 g90733(.A (n_8037), .B (n_2735), .C (csr_mcycle[21]), .D
       (n_2755), .E (csr_minstret[21]), .F (n_2733), .Q (n_2996));
  AN222X1 g90734(.A (n_2755), .B (csr_mcycle[9]), .C (csr_minstret[9]),
       .D (n_2733), .E (csr_mtvec[9]), .F (n_2731), .Q (n_2995));
  AO222X1 g90735(.A (csr_mcycle[39]), .B (n_2756), .C
       (csr_mscratch[7]), .D (n_2727), .E (csr_minstret[39]), .F
       (n_2732), .Q (n_2994));
  AO222X1 g90736(.A (n_8028), .B (n_2735), .C (csr_mcycle[11]), .D
       (n_2755), .E (csr_minstret[11]), .F (n_2733), .Q (n_2993));
  AO222X1 g90737(.A (csr_mtval[7]), .B (n_2726), .C (csr_mcycle[7]), .D
       (n_2755), .E (n_6256), .F (n_7370), .Q (n_2992));
  AO222X1 g90738(.A (n_8041), .B (n_2735), .C (csr_mcycle[24]), .D
       (n_2755), .E (csr_minstret[24]), .F (n_2733), .Q (n_2991));
  AN222X1 g90739(.A (n_2735), .B (n_8040), .C (csr_mcycle[55]), .D
       (n_2756), .E (csr_minstret[55]), .F (n_2732), .Q (n_2990));
  AO222X1 g90740(.A (n_8035), .B (n_2735), .C (csr_mcycle[19]), .D
       (n_2755), .E (csr_minstret[19]), .F (n_2733), .Q (n_2989));
  AO222X1 g90741(.A (n_8036), .B (n_2735), .C (csr_mcycle[20]), .D
       (n_2755), .E (csr_minstret[20]), .F (n_2733), .Q (n_2988));
  AN222X1 g90742(.A (n_2735), .B (n_8034), .C (csr_mcycle[18]), .D
       (n_2755), .E (csr_minstret[18]), .F (n_2733), .Q (n_2987));
  NA2X1 g90743(.A (n_2921), .B (n_2816), .Q (n_2986));
  AN222X1 g90744(.A (n_2755), .B (csr_mcycle[8]), .C (csr_minstret[8]),
       .D (n_2733), .E (csr_mtvec[8]), .F (n_2731), .Q (n_2985));
  NA2X1 g90745(.A (n_2944), .B (n_2861), .Q (n_2984));
  AO222X1 g90746(.A (n_8033), .B (n_2735), .C (csr_mcycle[49]), .D
       (n_2756), .E (csr_minstret[49]), .F (n_2732), .Q (n_2983));
  AO222X1 g90747(.A (n_8031), .B (n_2735), .C (csr_mcycle[16]), .D
       (n_2755), .E (csr_minstret[16]), .F (n_2733), .Q (n_2982));
  AN222X1 g90748(.A (n_2755), .B (csr_mcycle[6]), .C (csr_minstret[6]),
       .D (n_2733), .E (csr_mtvec[6]), .F (n_2731), .Q (n_2981));
  AN222X1 g90749(.A (n_2726), .B (csr_mtval[2]), .C (csr_mcycle[34]),
       .D (n_2756), .E (csr_minstret[34]), .F (n_2732), .Q (n_2980));
  AN221X1 g90750(.A (csr_minstret[3]), .B (n_2733), .C (csr_mtvec[3]),
       .D (n_2731), .E (n_2813), .Q (n_2979));
  AN222X1 g90751(.A (n_2755), .B (csr_mcycle[2]), .C (csr_minstret[2]),
       .D (n_2733), .E (csr_mtvec[2]), .F (n_2731), .Q (n_2978));
  AN222X1 g90752(.A (n_2756), .B (csr_mcycle[37]), .C
       (csr_minstret[37]), .D (n_2732), .E (n_7893), .F (n_2323), .Q
       (n_2977));
  AN222X1 g90754(.A (n_2756), .B (csr_mcycle[32]), .C
       (csr_minstret[32]), .D (n_2732), .E (csr_mtval[0]), .F (n_2726),
       .Q (n_2975));
  AN222X1 g90756(.A (n_2755), .B (csr_mcycle[5]), .C (csr_minstret[5]),
       .D (n_2733), .E (csr_mtvec[5]), .F (n_2731), .Q (n_2973));
  AN222X1 g90757(.A (n_2755), .B (csr_mcycle[4]), .C (csr_minstret[4]),
       .D (n_2733), .E (csr_mtvec[4]), .F (n_2731), .Q (n_2972));
  AN222X1 g90758(.A (n_2755), .B (csr_mcycle[0]), .C (csr_minstret[0]),
       .D (n_2733), .E (n_8051), .F (n_2731), .Q (n_2971));
  AN211X1 g90759(.A (n_2483), .B (n_2418), .C (n_2742), .D (n_2811), .Q
       (n_2970));
  NO3X1 g90760(.A (n_2859), .B (n_2920), .C (n_2307), .Q (n_3006));
  NO2X4 g90761(.A (n_2331), .B (n_2304), .Q (n_2334));
  NO2X4 g90762(.A (n_8659), .B (n_2305), .Q (n_2333));
  NO2X4 g90763(.A (n_2331), .B (n_2305), .Q (n_3004));
  NO2X4 g90764(.A (n_8659), .B (n_2304), .Q (n_2332));
  INX1 g90765(.A (n_2969), .Q (n_2968));
  AN221X1 g90766(.A (csr_mscratch[19]), .B (n_2727), .C (n_7907), .D
       (n_2323), .E (n_2868), .Q (n_2967));
  AN22X1 g90767(.A (n_2756), .B (csr_mcycle[59]), .C (n_2732), .D
       (csr_minstret[59]), .Q (n_2966));
  AN22X1 g90768(.A (n_2756), .B (csr_mcycle[61]), .C (n_2732), .D
       (csr_minstret[61]), .Q (n_2965));
  NO2X1 g90769(.A (n_957), .B (n_7714), .Q (n_2964));
  AN221X1 g90770(.A (csr_mscratch[5]), .B (n_2727), .C (csr_mtval[5]),
       .D (n_2726), .E (n_2821), .Q (n_2963));
  AN221X1 g90771(.A (csr_mscratch[6]), .B (n_2727), .C (csr_mtval[6]),
       .D (n_2726), .E (n_2834), .Q (n_2962));
  AN221X1 g90773(.A (csr_mcause[22]), .B (n_2725), .C (csr_mtval[22]),
       .D (n_2726), .E (n_2883), .Q (n_2960));
  AN221X1 g90774(.A (csr_mcause[26]), .B (n_2725), .C (csr_mtval[26]),
       .D (n_2726), .E (n_2881), .Q (n_2959));
  AN221X1 g90775(.A (csr_mscratch[31]), .B (n_2727), .C (n_7911), .D
       (n_2323), .E (n_2878), .Q (n_2958));
  AN221X1 g90776(.A (csr_mcause[11]), .B (n_2725), .C (csr_mtval[11]),
       .D (n_2726), .E (n_2869), .Q (n_2957));
  AN221X1 g90777(.A (csr_mscratch[24]), .B (n_2727), .C (n_7885), .D
       (n_2323), .E (n_2866), .Q (n_2956));
  AN221X1 g90778(.A (csr_mscratch[9]), .B (n_2727), .C (csr_mtval[9]),
       .D (n_2726), .E (n_2842), .Q (n_2955));
  AN221X1 g90779(.A (csr_mscratch[21]), .B (n_2727), .C (n_7909), .D
       (n_2323), .E (n_2867), .Q (n_2954));
  AN221X1 g90780(.A (csr_mscratch[14]), .B (n_2727), .C
       (csr_mtval[14]), .D (n_2726), .E (n_2847), .Q (n_2953));
  AN221X1 g90781(.A (csr_mcause[13]), .B (n_2725), .C (n_7901), .D
       (n_2323), .E (n_2845), .Q (n_2952));
  AN221X1 g90782(.A (csr_mcause[15]), .B (n_2725), .C (n_7903), .D
       (n_2323), .E (n_2846), .Q (n_2951));
  AN221X1 g90783(.A (csr_mcause[16]), .B (n_2725), .C (csr_mtval[16]),
       .D (n_2726), .E (n_2824), .Q (n_2950));
  AN221X1 g90784(.A (csr_mcause[20]), .B (n_2725), .C (csr_mtval[20]),
       .D (n_2726), .E (n_2864), .Q (n_2949));
  AN221X1 g90785(.A (csr_mscratch[10]), .B (n_2727), .C
       (csr_mtval[10]), .D (n_2726), .E (n_2844), .Q (n_2948));
  NA2X2 g90786(.A (n_8566), .B (n_7282), .Q (n_7707));
  NA2X2 g90787(.A (n_8566), .B (n_958), .Q (n_7708));
  OR2X2 g90788(.A (n_8566), .B (n_958), .Q (n_7710));
  NO2X2 g90789(.A (n_8566), .B (n_7282), .Q (n_8165));
  NA2X1 g90790(.A (n_8566), .B (n_2635), .Q (n_2969));
  INX1 g90791(.A (n_2946), .Q (n_2947));
  INX2 g90792(.A (n_2942), .Q (n_2943));
  INX3 g90795(.A (n_2938), .Q (n_2937));
  AN22X1 g90797(.A (n_2756), .B (csr_mcycle[62]), .C (n_2732), .D
       (csr_minstret[62]), .Q (n_2934));
  AN22X1 g90798(.A (n_2756), .B (csr_mcycle[57]), .C (n_2732), .D
       (csr_minstret[57]), .Q (n_2933));
  AN22X1 g90799(.A (n_2756), .B (csr_mcycle[50]), .C (n_2732), .D
       (csr_minstret[50]), .Q (n_2932));
  ON21X1 g90800(.A (n_2728), .B (n_6084), .C (n_2817), .Q (n_2931));
  AN22X1 g90801(.A (n_2755), .B (csr_mcycle[17]), .C (n_2733), .D
       (csr_minstret[17]), .Q (n_2930));
  AN22X1 g90802(.A (n_2755), .B (csr_mcycle[23]), .C (n_2733), .D
       (csr_minstret[23]), .Q (n_2929));
  AN221X1 g90803(.A (csr_minstret[7]), .B (n_2733), .C (csr_mtvec[7]),
       .D (n_2731), .E (n_2768), .Q (n_2928));
  AN22X1 g90804(.A (n_2756), .B (csr_mcycle[40]), .C (n_2732), .D
       (csr_minstret[40]), .Q (n_2927));
  AN221X1 g90805(.A (csr_utime[1]), .B (n_2619), .C (csr_mcause[1]), .D
       (n_2725), .E (n_2766), .Q (n_2926));
  AND3X1 g90806(.A (n_2812), .B (n_2694), .C (n_2693), .Q (n_2925));
  AN22X1 g90807(.A (n_2756), .B (csr_mcycle[33]), .C (n_2732), .D
       (csr_minstret[33]), .Q (n_2924));
  AN22X1 g90809(.A (n_2756), .B (csr_mcycle[60]), .C (n_2732), .D
       (csr_minstret[60]), .Q (n_2922));
  AN22X1 g90810(.A (n_2756), .B (csr_mcycle[36]), .C (n_2732), .D
       (csr_minstret[36]), .Q (n_2921));
  NO2X1 g90811(.A (n_2329), .B (n_8157), .Q (n_2920));
  OR5X1 g90812(.A (n_2329), .B (n_2577), .C (store_type), .D
       (branch_type), .E (system_type), .Q (n_2919));
  NA3I1X1 g90813(.B (n_2858), .C (n_2703), .AN (n_2696), .Q (n_2918));
  NO2I1X1 g90814(.B (n_2701), .AN (n_2860), .Q (n_2946));
  NA2I1X1 g90815(.B (n_8569), .AN (n_2859), .Q (n_2945));
  AND2X1 g90816(.A (n_2858), .B (n_2763), .Q (n_2944));
  NO2I1X4 g90817(.B (n_2330), .AN (n_2852), .Q (n_2942));
  NO2X4 g90819(.A (n_2330), .B (n_2851), .Q (n_2939));
  AND2X4 g90820(.A (n_2757), .B (n_2855), .Q (n_2938));
  NO2X4 g90821(.A (n_2330), .B (n_2857), .Q (n_2936));
  INX2 g90824(.A (n_2330), .Q (n_2917));
  INX8 g90825(.A (n_2757), .Q (n_2330));
  INX1 g90826(.A (n_2916), .Q (n_7272));
  INX1 g90827(.A (n_2915), .Q (n_7273));
  INX1 g90828(.A (n_2914), .Q (n_7278));
  INX1 g90829(.A (n_2913), .Q (n_7263));
  INX1 g90830(.A (n_2912), .Q (n_7280));
  INX1 g90831(.A (n_2911), .Q (n_7279));
  INX1 g90832(.A (n_2910), .Q (n_7257));
  INX1 g90833(.A (n_2909), .Q (n_7264));
  INX1 g90834(.A (n_2908), .Q (n_7261));
  INX2 g90835(.A (n_2907), .Q (n_7251));
  INX1 g90836(.A (n_2906), .Q (n_7250));
  INX1 g90837(.A (n_2905), .Q (n_7252));
  INX1 g90838(.A (n_2904), .Q (n_7253));
  INX1 g90839(.A (n_2903), .Q (n_7254));
  INX1 g90840(.A (n_2902), .Q (n_7255));
  INX1 g90841(.A (n_2901), .Q (n_7256));
  INX1 g90842(.A (n_2900), .Q (n_7258));
  INX1 g90843(.A (n_2899), .Q (n_7259));
  INX1 g90844(.A (n_2898), .Q (n_7260));
  INX1 g90845(.A (n_2897), .Q (n_7262));
  INX1 g90846(.A (n_2896), .Q (n_7265));
  INX1 g90847(.A (n_2895), .Q (n_7270));
  INX1 g90848(.A (n_2894), .Q (n_7271));
  INX1 g90849(.A (n_2893), .Q (n_7274));
  INX1 g90850(.A (n_2892), .Q (n_7267));
  INX1 g90851(.A (n_2891), .Q (n_7277));
  INX1 g90852(.A (n_2890), .Q (n_7268));
  INX1 g90853(.A (n_2889), .Q (n_7269));
  INX1 g90854(.A (n_2888), .Q (n_7266));
  INX1 g90855(.A (n_2887), .Q (n_7276));
  INX1 g90856(.A (n_958), .Q (n_7282));
  AN22X1 g90858(.A (n_2727), .B (csr_mscratch[27]), .C (n_2323), .D
       (n_7888), .Q (n_2885));
  AN22X1 g90859(.A (n_2727), .B (csr_mscratch[17]), .C (n_2323), .D
       (n_7905), .Q (n_2884));
  AO22X1 g90860(.A (n_2727), .B (csr_mscratch[22]), .C (n_2323), .D
       (n_7910), .Q (n_2883));
  AN22X1 g90861(.A (n_2727), .B (csr_mscratch[30]), .C (n_2323), .D
       (n_7900), .Q (n_2882));
  AO22X1 g90862(.A (n_2727), .B (csr_mscratch[26]), .C (n_2323), .D
       (n_7887), .Q (n_2881));
  AN22X1 g90863(.A (n_2725), .B (csr_mcause[30]), .C (n_2726), .D
       (csr_mtval[30]), .Q (n_2880));
  AN22X1 g90864(.A (n_2725), .B (csr_mcause[28]), .C (n_2726), .D
       (csr_mtval[28]), .Q (n_2879));
  AO22X1 g90865(.A (n_2725), .B (csr_mcause[31]), .C (n_2726), .D
       (csr_mtval[31]), .Q (n_2878));
  AN22X1 g90866(.A (n_2725), .B (csr_mcause[29]), .C (n_2726), .D
       (csr_mtval[29]), .Q (n_2877));
  AN22X1 g90867(.A (n_2727), .B (csr_mscratch[29]), .C (n_2323), .D
       (n_7891), .Q (n_2876));
  AN22X1 g90868(.A (n_2727), .B (csr_mscratch[28]), .C (n_2323), .D
       (n_7889), .Q (n_2875));
  AN22X1 g90869(.A (n_2725), .B (csr_mcause[27]), .C (n_2726), .D
       (csr_mtval[27]), .Q (n_2874));
  AN22X1 g90870(.A (n_2725), .B (csr_mcause[23]), .C (n_2726), .D
       (csr_mtval[23]), .Q (n_2873));
  AN22X1 g90871(.A (n_2725), .B (csr_mcause[25]), .C (n_2726), .D
       (csr_mtval[25]), .Q (n_2872));
  AO22X1 g90872(.A (n_2725), .B (csr_mcause[12]), .C (n_2323), .D
       (n_7899), .Q (n_2871));
  AN22X1 g90873(.A (n_2727), .B (csr_mscratch[25]), .C (n_2323), .D
       (n_7886), .Q (n_2870));
  AO22X1 g90874(.A (n_2727), .B (csr_mscratch[11]), .C (n_2323), .D
       (n_7898), .Q (n_2869));
  AO22X1 g90875(.A (n_2725), .B (csr_mcause[19]), .C (n_2726), .D
       (csr_mtval[19]), .Q (n_2868));
  AO22X1 g90876(.A (n_2725), .B (csr_mcause[21]), .C (n_2726), .D
       (csr_mtval[21]), .Q (n_2867));
  AO22X1 g90877(.A (n_2725), .B (csr_mcause[24]), .C (n_2726), .D
       (csr_mtval[24]), .Q (n_2866));
  ON21X1 g90878(.A (n_2728), .B (n_2484), .C (n_2503), .Q (n_8177));
  AN22X1 g90879(.A (n_2727), .B (csr_mscratch[23]), .C (n_2323), .D
       (n_7884), .Q (n_2865));
  AO22X1 g90880(.A (n_2727), .B (csr_mscratch[20]), .C (n_2323), .D
       (n_7908), .Q (n_2864));
  AN22X1 g90881(.A (n_2727), .B (csr_mscratch[18]), .C (n_2323), .D
       (n_7906), .Q (n_2863));
  AN22X1 g90882(.A (n_2725), .B (csr_mcause[17]), .C (n_2726), .D
       (csr_mtval[17]), .Q (n_2862));
  MU2IX1 g90883(.S (n_2722), .IN0 (n_7816), .IN1 (n_7815), .Q (n_2916));
  MU2IX1 g90884(.S (n_2722), .IN0 (n_7818), .IN1 (n_7817), .Q (n_2915));
  MU2IX1 g90885(.S (n_2722), .IN0 (n_7820), .IN1 (n_7819), .Q (n_2914));
  MU2IX1 g90886(.S (n_2322), .IN0 (n_7792), .IN1 (n_7791), .Q (n_2913));
  MU2IX1 g90887(.S (n_2722), .IN0 (n_7824), .IN1 (n_7823), .Q (n_2912));
  MU2IX1 g90888(.S (n_2722), .IN0 (n_7822), .IN1 (n_7821), .Q (n_2911));
  MU2IX1 g90889(.S (n_2322), .IN0 (n_7780), .IN1 (n_7779), .Q (n_2910));
  MU2IX1 g90890(.S (n_2322), .IN0 (n_7794), .IN1 (n_7793), .Q (n_2909));
  MU2IX1 g90891(.S (n_2322), .IN0 (n_7788), .IN1 (n_7787), .Q (n_2908));
  MU2IX1 g90892(.S (n_2322), .IN0 (n_7766), .IN1 (n_7765), .Q (n_2907));
  MU2IX1 g90893(.S (n_2322), .IN0 (n_7768), .IN1 (n_7767), .Q (n_2906));
  MU2IX1 g90894(.S (n_2322), .IN0 (n_7770), .IN1 (n_7769), .Q (n_2905));
  MU2IX1 g90895(.S (n_2322), .IN0 (n_7772), .IN1 (n_7771), .Q (n_2904));
  MU2IX1 g90896(.S (n_2322), .IN0 (n_7774), .IN1 (n_7773), .Q (n_2903));
  MU2IX1 g90897(.S (n_2322), .IN0 (n_7776), .IN1 (n_7775), .Q (n_2902));
  MU2IX1 g90898(.S (n_2322), .IN0 (n_7778), .IN1 (n_7777), .Q (n_2901));
  MU2IX1 g90899(.S (n_2322), .IN0 (n_7782), .IN1 (n_7781), .Q (n_2900));
  MU2IX1 g90900(.S (n_2322), .IN0 (n_7784), .IN1 (n_7783), .Q (n_2899));
  MU2IX1 g90901(.S (n_2322), .IN0 (n_7786), .IN1 (n_7785), .Q (n_2898));
  MU2IX1 g90902(.S (n_2322), .IN0 (n_7790), .IN1 (n_7789), .Q (n_2897));
  MU2IX1 g90903(.S (n_2322), .IN0 (n_7796), .IN1 (n_7795), .Q (n_2896));
  MU2IX1 g90904(.S (n_2722), .IN0 (n_7808), .IN1 (n_7807), .Q (n_2895));
  MU2IX1 g90905(.S (n_2322), .IN0 (n_7810), .IN1 (n_7809), .Q (n_2894));
  MU2IX1 g90906(.S (n_2322), .IN0 (n_7806), .IN1 (n_7805), .Q (n_2893));
  MU2IX1 g90907(.S (n_2322), .IN0 (n_7798), .IN1 (n_7797), .Q (n_2892));
  MU2IX1 g90908(.S (n_2322), .IN0 (n_7804), .IN1 (n_7803), .Q (n_2891));
  MU2IX1 g90909(.S (n_2322), .IN0 (n_7800), .IN1 (n_7799), .Q (n_2890));
  MU2IX1 g90910(.S (n_2322), .IN0 (n_7802), .IN1 (n_7801), .Q (n_2889));
  MU2IX1 g90911(.S (n_2322), .IN0 (n_7812), .IN1 (n_7811), .Q (n_2888));
  MU2IX1 g90912(.S (n_2322), .IN0 (n_7814), .IN1 (n_7813), .Q (n_2887));
  MU2IX2 g90913(.S (n_2721), .IN0 (n_7828), .IN1 (n_7827), .Q (n_958));
  INX2 g90917(.A (n_2855), .Q (n_2856));
  INX1 g90918(.A (n_2853), .Q (n_2854));
  INX2 g90919(.A (n_2852), .Q (n_2853));
  INX1 g90920(.A (n_2851), .Q (n_2850));
  INX4 g90942(.A (n_2326), .Q (alu_operation_code_39112));
  AO221X1 g90943(.A (csr_utime[12]), .B (n_2619), .C (n_2313), .D
       (csr_utime[44]), .E (n_7370), .Q (n_2849));
  AN22X1 g90944(.A (n_2725), .B (csr_mcause[18]), .C (n_2726), .D
       (csr_mtval[18]), .Q (n_2848));
  AO222X1 g90945(.A (csr_utime[14]), .B (n_2619), .C (csr_mcause[14]),
       .D (n_2725), .E (csr_utime[46]), .F (n_2312), .Q (n_2847));
  ON221X1 g90946(.A (n_2484), .B (n_2724), .C (n_7714), .D (n_8078), .E
       (n_2503), .Q (n_8205));
  AO222X1 g90947(.A (csr_utime[15]), .B (n_2619), .C
       (csr_mscratch[15]), .D (n_2727), .E (csr_utime[47]), .F
       (n_2312), .Q (n_2846));
  AO222X1 g90948(.A (csr_utime[13]), .B (n_2619), .C
       (csr_mscratch[13]), .D (n_2727), .E (csr_utime[45]), .F
       (n_2313), .Q (n_2845));
  AO222X1 g90949(.A (csr_utime[10]), .B (n_2619), .C (csr_mcause[10]),
       .D (n_2725), .E (csr_utime[42]), .F (n_2313), .Q (n_2844));
  ON21X1 g90950(.A (n_2325), .B (n_4442), .C (n_2775), .Q (n_2843));
  AO222X1 g90951(.A (csr_utime[9]), .B (n_2619), .C (csr_mcause[9]), .D
       (n_2725), .E (csr_utime[41]), .F (n_2312), .Q (n_2842));
  AN22X1 g90952(.A (n_2725), .B (csr_mcause[8]), .C (n_2726), .D
       (csr_mtval[8]), .Q (n_2841));
  AO222X1 g90953(.A (csr_utime[26]), .B (n_2619), .C (n_4446), .D
       (n_2324), .E (csr_utime[58]), .F (n_2313), .Q (n_2840));
  AN222X1 g90954(.A (n_2619), .B (csr_utime[28]), .C (csr_utime[60]),
       .D (n_2313), .E (n_4448), .F (n_2324), .Q (n_2839));
  ON21X1 g90955(.A (n_8358), .B (n_2484), .C (n_2503), .Q (n_8170));
  ON222X1 g90956(.A (csr_utime[31]), .B (n_2620), .C (n_4451), .D
       (n_2325), .E (n_2314), .F (csr_utime[63]), .Q (n_2838));
  AN222X1 g90957(.A (n_2619), .B (csr_utime[29]), .C (csr_utime[61]),
       .D (n_2614), .E (n_4449), .F (n_2324), .Q (n_2837));
  AN222X1 g90958(.A (n_2619), .B (csr_utime[27]), .C (csr_utime[59]),
       .D (n_2313), .E (n_4447), .F (n_2324), .Q (n_2836));
  AN222X1 g90959(.A (n_2619), .B (csr_utime[25]), .C (csr_utime[57]),
       .D (n_2313), .E (n_4445), .F (n_2324), .Q (n_2835));
  AO222X1 g90960(.A (csr_utime[6]), .B (n_2619), .C (csr_mcause[6]), .D
       (n_2725), .E (csr_utime[38]), .F (n_2312), .Q (n_2834));
  ON222X1 g90961(.A (csr_utime[21]), .B (n_2620), .C (n_4441), .D
       (n_2325), .E (n_2615), .F (csr_utime[53]), .Q (n_2833));
  AN222X1 g90962(.A (n_2619), .B (csr_utime[23]), .C (csr_utime[55]),
       .D (n_2313), .E (n_4443), .F (n_2324), .Q (n_2832));
  ON222X1 g90963(.A (csr_utime[20]), .B (n_2620), .C (n_4440), .D
       (n_2325), .E (n_2615), .F (csr_utime[52]), .Q (n_2831));
  AN222X1 g90964(.A (n_2619), .B (csr_utime[18]), .C (csr_utime[50]),
       .D (n_2312), .E (n_4438), .F (n_2324), .Q (n_2830));
  ON222X1 g90965(.A (csr_utime[24]), .B (n_2620), .C (n_4444), .D
       (n_2325), .E (n_2615), .F (csr_utime[56]), .Q (n_2829));
  ON222X1 g90966(.A (csr_utime[19]), .B (n_2620), .C (n_4439), .D
       (n_2325), .E (n_2314), .F (csr_utime[51]), .Q (n_2828));
  ON21X1 g90967(.A (n_2734), .B (n_2484), .C (n_2503), .Q (n_8169));
  AN222X1 g90968(.A (n_2619), .B (csr_utime[17]), .C (csr_utime[49]),
       .D (n_2313), .E (n_4437), .F (n_2324), .Q (n_2827));
  ON222X1 g90969(.A (csr_utime[16]), .B (n_2620), .C (n_4436), .D
       (n_2325), .E (n_2314), .F (csr_utime[48]), .Q (n_2826));
  AN221X1 g90970(.A (csr_utime[62]), .B (n_2614), .C (csr_utime[30]),
       .D (n_2619), .E (n_2744), .Q (n_2825));
  AO22X1 g90971(.A (n_2727), .B (csr_mscratch[16]), .C (n_2323), .D
       (n_7904), .Q (n_2824));
  AN22X1 g90972(.A (n_2725), .B (csr_mcause[4]), .C (n_2726), .D
       (csr_mtval[4]), .Q (n_2823));
  ON221X1 g90973(.A (csr_utime[11]), .B (n_2620), .C (csr_utime[43]),
       .D (n_2314), .E (n_2736), .Q (n_2822));
  AO222X1 g90974(.A (csr_utime[5]), .B (n_2619), .C (csr_mcause[5]), .D
       (n_2725), .E (csr_utime[37]), .F (n_2313), .Q (n_2821));
  AO21X1 g90975(.A (n_2732), .B (csr_minstret[35]), .C (n_2747), .Q
       (n_2820));
  AN221X1 g90976(.A (csr_utime[40]), .B (n_2313), .C (csr_utime[8]), .D
       (n_2619), .E (n_2744), .Q (n_2819));
  AO22X1 g90977(.A (n_2324), .B (n_4435), .C (n_2735), .D (n_8030), .Q
       (n_2818));
  AN21X1 g90978(.A (n_2619), .B (csr_utime[2]), .C (n_2767), .Q
       (n_2817));
  AN221X1 g90979(.A (csr_utime[36]), .B (n_2614), .C (csr_utime[4]), .D
       (n_2619), .E (n_2738), .Q (n_2816));
  AND2X1 g90980(.A (n_2758), .B (n_2596), .Q (n_2815));
  NA3X1 g90981(.A (n_2699), .B (n_2691), .C (n_7882), .Q (n_2814));
  AO22X1 g90982(.A (n_7370), .B (n_7275), .C (n_2619), .D
       (csr_utime[3]), .Q (n_2813));
  NO3I1X1 g90983(.B (n_2707), .C (n_2709), .AN (n_2700), .Q (n_2812));
  AO222X1 g90984(.A (store_type), .B (n_2514), .C (n_2497), .D
       (n_2712), .E (n_2308), .F (branch_type), .Q (n_2811));
  NA3X1 g90985(.A (n_2707), .B (n_2694), .C (n_2693), .Q (n_2810));
  NO3I1X1 g90986(.B (n_2699), .C (n_2705), .AN (n_2691), .Q (n_2809));
  NA3I1X1 g90987(.B (n_2760), .C (n_7275), .AN (n_2700), .Q (n_2808));
  NA3I2X1 g90988(.C (n_2692), .AN (n_2759), .BN (n_2697), .Q (n_2807));
  AND2X1 g90990(.A (n_2762), .B (n_2765), .Q (n_2861));
  NO3I1X1 g90992(.B (n_2699), .C (n_2698), .AN (n_2691), .Q (n_2860));
  AN21X1 g90993(.A (prev_load_request), .B (read_response), .C
       (n_2758), .Q (n_2859));
  NO3I2X1 g90994(.C (n_2759), .AN (n_2697), .BN (n_2692), .Q (n_2858));
  OR2X4 g90995(.A (n_2684), .B (n_2510), .Q (n_2857));
  NO2X4 g90996(.A (n_2803), .B (n_2510), .Q (n_2855));
  NO2I1X4 g90997(.B (n_2803), .AN (n_2510), .Q (n_2852));
  NA2X4 g90998(.A (n_2803), .B (n_2510), .Q (n_2851));
  NA2X4 g90999(.A (n_2764), .B (n_8484), .Q (n_2326));
  INX1 g91000(.A (n_2805), .Q (n_2804));
  INX4 g91001(.A (n_2684), .Q (n_2803));
  HAX1 g91002(.A (n_2488), .B (n_2441), .S (n_2805), .CO (n_2802));
  AO222X1 g91003(.A (csr_mtvec[14]), .B (n_2569), .C (n_2568), .D
       (n_7846), .E (n_960), .F (n_7902), .Q (n_2801));
  AO222X1 g91005(.A (csr_mtvec[27]), .B (n_2569), .C (n_2568), .D
       (n_7833), .E (n_960), .F (n_7888), .Q (n_2799));
  AO222X1 g91006(.A (csr_mtvec[23]), .B (n_2569), .C (n_2568), .D
       (n_7837), .E (n_960), .F (n_7884), .Q (n_2798));
  AO222X1 g91007(.A (csr_mtvec[19]), .B (n_2569), .C (n_2568), .D
       (n_7841), .E (n_960), .F (n_7907), .Q (n_2797));
  AO222X1 g91008(.A (csr_mtvec[31]), .B (n_2569), .C (n_2568), .D
       (n_7829), .E (n_960), .F (n_7911), .Q (n_2796));
  AO222X1 g91009(.A (csr_mtvec[30]), .B (n_2569), .C (n_2568), .D
       (n_7830), .E (n_960), .F (n_7900), .Q (n_2795));
  AO222X1 g91010(.A (csr_mtvec[29]), .B (n_2569), .C (n_2568), .D
       (n_7831), .E (n_960), .F (n_7891), .Q (n_2794));
  AO222X1 g91011(.A (csr_mtvec[26]), .B (n_2569), .C (n_2568), .D
       (n_7834), .E (n_960), .F (n_7887), .Q (n_2793));
  AO222X1 g91012(.A (csr_mtvec[25]), .B (n_2569), .C (n_2568), .D
       (n_7835), .E (n_960), .F (n_7886), .Q (n_2792));
  AO222X1 g91013(.A (csr_mtvec[22]), .B (n_2569), .C (n_2568), .D
       (n_7838), .E (n_960), .F (n_7910), .Q (n_2791));
  AO222X1 g91014(.A (csr_mtvec[21]), .B (n_2569), .C (n_2568), .D
       (n_7839), .E (n_960), .F (n_7909), .Q (n_2790));
  AO222X1 g91015(.A (csr_mtvec[18]), .B (n_2569), .C (n_2568), .D
       (n_7842), .E (n_960), .F (n_7906), .Q (n_2789));
  AO222X1 g91016(.A (csr_mtvec[15]), .B (n_2569), .C (n_2568), .D
       (n_7845), .E (n_960), .F (n_7903), .Q (n_2788));
  AO222X1 g91017(.A (csr_mtvec[28]), .B (n_2569), .C (n_2568), .D
       (n_7832), .E (n_960), .F (n_7889), .Q (n_2787));
  AO222X1 g91018(.A (csr_mtvec[24]), .B (n_2569), .C (n_2568), .D
       (n_7836), .E (n_960), .F (n_7885), .Q (n_2786));
  AO222X1 g91019(.A (csr_mtvec[20]), .B (n_2569), .C (n_2568), .D
       (n_7840), .E (n_960), .F (n_7908), .Q (n_2785));
  AO222X1 g91020(.A (csr_mtvec[17]), .B (n_2569), .C (n_2568), .D
       (n_7843), .E (n_960), .F (n_7905), .Q (n_2784));
  AO222X1 g91022(.A (csr_mtvec[11]), .B (n_2569), .C (n_2568), .D
       (n_7849), .E (n_960), .F (n_7898), .Q (n_2782));
  AO222X1 g91023(.A (csr_mtvec[16]), .B (n_2569), .C (n_2568), .D
       (n_7844), .E (n_960), .F (n_7904), .Q (n_2781));
  NA2I1X1 g91024(.B (n_2323), .AN (n_2484), .Q (n_2780));
  NA2I1X0 g91025(.B (n_2726), .AN (n_2484), .Q (n_2779));
  AO222X1 g91026(.A (csr_mtvec[13]), .B (n_2569), .C (n_2568), .D
       (n_7847), .E (n_960), .F (n_7901), .Q (n_2778));
  AO222X1 g91027(.A (csr_mtvec[10]), .B (n_2569), .C (n_2568), .D
       (n_7850), .E (n_960), .F (n_7897), .Q (n_2777));
  NA2X1 g91028(.A (n_2731), .B (csr_mtvec[25]), .Q (n_2776));
  AN22X1 g91029(.A (n_2619), .B (csr_utime[22]), .C (n_2313), .D
       (csr_utime[54]), .Q (n_2775));
  NA2X1 g91030(.A (n_2731), .B (csr_mtvec[23]), .Q (n_2774));
  NA2X1 g91031(.A (n_2731), .B (csr_mtvec[18]), .Q (n_2773));
  AO222X1 g91032(.A (csr_mtvec[12]), .B (n_2569), .C (n_2568), .D
       (n_7848), .E (n_960), .F (n_7899), .Q (n_2772));
  AO222X1 g91033(.A (csr_mtvec[9]), .B (n_2569), .C (n_2568), .D
       (n_7851), .E (n_960), .F (n_7896), .Q (n_2771));
  ON22X1 g91036(.A (n_2620), .B (csr_utime[7]), .C (n_2314), .D
       (csr_utime[39]), .Q (n_2768));
  ON21X1 g91037(.A (n_2314), .B (csr_utime[34]), .C (n_2741), .Q
       (n_2767));
  ON21X1 g91038(.A (n_2314), .B (csr_utime[33]), .C (n_2741), .Q
       (n_2766));
  INX1 g91039(.A (n_2761), .Q (n_2762));
  INX8 g91040(.A (n_2746), .Q (n_2756));
  INX8 g91041(.A (n_2745), .Q (n_2755));
  NO2X2 g91042(.A (n_2687), .B (n_2480), .Q (irq_fast_response[11]));
  AO222X1 g91043(.A (csr_mtvec[8]), .B (n_2569), .C (n_2568), .D
       (n_7852), .E (n_960), .F (n_7895), .Q (n_2754));
  NO2X2 g91044(.A (n_2689), .B (n_2480), .Q (irq_fast_response[15]));
  AO222X1 g91045(.A (csr_mtvec[7]), .B (n_2569), .C (n_2568), .D
       (n_7853), .E (n_960), .F (n_7923), .Q (n_2753));
  AND2X1 g91046(.A (n_2690), .B (n_2486), .Q (irq_fast_response[13]));
  AND2X1 g91047(.A (n_2690), .B (n_2485), .Q (irq_fast_response[14]));
  AND2X1 g91048(.A (n_2686), .B (n_2486), .Q (irq_fast_response[5]));
  AND2X1 g91051(.A (n_2686), .B (n_2485), .Q (irq_fast_response[6]));
  AO222X1 g91052(.A (csr_mtvec[6]), .B (n_2569), .C (n_2568), .D
       (n_7854), .E (n_960), .F (n_7894), .Q (n_2752));
  AO222X1 g91053(.A (csr_mtvec[5]), .B (n_2569), .C (n_2568), .D
       (n_7855), .E (n_960), .F (n_7893), .Q (n_2751));
  AO222X1 g91054(.A (csr_mtvec[4]), .B (n_2569), .C (n_2568), .D
       (n_7856), .E (n_960), .F (n_7892), .Q (n_2750));
  AO222X1 g91055(.A (csr_mtvec[3]), .B (n_2569), .C (n_2568), .D
       (n_7857), .E (n_960), .F (n_7964), .Q (n_2749));
  AO222X1 g91056(.A (n_8664), .B (n_2568), .C (csr_mtvec[2]), .D
       (n_2569), .E (n_960), .F (n_7890), .Q (n_2748));
  AND2X1 g91057(.A (n_2688), .B (n_2485), .Q (irq_fast_response[10]));
  AND2X1 g91058(.A (n_2688), .B (n_2486), .Q (irq_fast_response[9]));
  AND2X1 g91059(.A (n_2688), .B (n_2482), .Q (irq_fast_response[8]));
  ON21X1 g91060(.A (n_2314), .B (csr_utime[35]), .C (n_2737), .Q
       (n_2747));
  AND2X1 g91061(.A (n_2685), .B (n_2479), .Q (irq_fast_response[3]));
  AND2X1 g91062(.A (n_2685), .B (n_2485), .Q (irq_fast_response[2]));
  AND2X1 g91063(.A (n_2685), .B (n_2486), .Q (irq_fast_response[1]));
  AND2X1 g91064(.A (n_2685), .B (n_2482), .Q (irq_fast_response[0]));
  AND2X1 g91065(.A (n_2690), .B (n_2482), .Q (irq_fast_response[12]));
  AND2X1 g91066(.A (n_2686), .B (n_2482), .Q (irq_fast_response[4]));
  AND2X1 g91067(.A (n_2686), .B (n_2479), .Q (irq_fast_response[7]));
  NA2I1X1 g91068(.B (n_7275), .AN (n_2702), .Q (n_2765));
  NA2X1 g91069(.A (n_2720), .B (n_2487), .Q (n_2764));
  NO2X1 g91070(.A (n_2703), .B (n_2696), .Q (n_2763));
  NO2I1X1 g91071(.B (n_2704), .AN (n_7275), .Q (n_2761));
  NA2I1X1 g91072(.B (n_7275), .AN (n_2706), .Q (n_2760));
  NA2X1 g91073(.A (n_2708), .B (n_2695), .Q (n_2759));
  OR2X1 g91074(.A (n_2742), .B (n_8073), .Q (n_2758));
  NA2I1X4 g91075(.B (n_2683), .AN (n_8164), .Q (n_2757));
  NA2X2 g91076(.A (n_2743), .B (n_2508), .Q (n_2746));
  NA2X4 g91077(.A (n_2743), .B (n_2591), .Q (n_2745));
  INX1 g91079(.A (n_2737), .Q (n_2738));
  INX1 g91080(.A (n_7370), .Q (n_2736));
  INX1 g91088(.A (n_2324), .Q (n_2325));
  INX4 g91089(.A (n_2734), .Q (n_2735));
  INX8 g91090(.A (n_2711), .Q (n_2733));
  INX4 g91091(.A (n_2710), .Q (n_2732));
  INX6 g91092(.A (n_8358), .Q (n_2731));
  BUX4 g91100(.A (n_2729), .Q (n_2323));
  INX8 g91101(.A (n_2728), .Q (n_2727));
  INX6 g91102(.A (n_2260), .Q (n_2726));
  INX4 g91103(.A (n_2724), .Q (n_2725));
  BUCX8 g91106(.A (n_2722), .Q (n_2322));
  INX1 g91107(.A (n_2321), .Q (n_2722));
  INX1 g91112(.A (n_2721), .Q (n_2321));
  OR5X1 g91113(.A (n_8159), .B (n_8158), .C (n_8161), .D (n_8163), .E
       (n_2308), .Q (n_2720));
  NA2X4 g91114(.A (n_2259), .B (n_2642), .Q (n_2719));
  AN21X1 g91115(.A (n_6121), .B (n_2589), .C (n_2641), .Q (n_2718));
  NO2X2 g91118(.A (n_2581), .B (n_2647), .Q (n_2715));
  NA2X2 g91119(.A (n_2654), .B (n_2644), .Q (n_2714));
  NA2X2 g91120(.A (n_2653), .B (n_2645), .Q (n_2713));
  NO2X1 g91121(.A (n_2638), .B (n_2509), .Q (n_7694));
  ON21X1 g91122(.A (n_2597), .B (n_8163), .C (n_2595), .Q (n_2712));
  NA2X1 g91123(.A (n_2637), .B (n_2591), .Q (n_3869_BAR));
  NO2X1 g91124(.A (n_2625), .B (n_2277), .Q (n_2744));
  NO2X2 g91125(.A (n_2600), .B (n_2622), .Q (n_2743));
  AN31X1 g91126(.A (n_2505), .B (n_2511), .C (n_8309), .D (n_8073), .Q
       (n_2742));
  NA2X1 g91127(.A (n_2636), .B (n_2599), .Q (n_2741));
  NO2X1 g91128(.A (n_2513), .B (n_2622), .Q (n_2739));
  NA2X1 g91129(.A (n_2636), .B (n_2592), .Q (n_2737));
  NO2X2 g91131(.A (n_2625), .B (n_2622), .Q (n_7370));
  NO2X4 g91132(.A (n_2623), .B (n_2634), .Q (n_2324));
  OR2X2 g91133(.A (n_2625), .B (n_2634), .Q (n_2734));
  NA2X4 g91134(.A (n_2631), .B (n_2591), .Q (n_2711));
  NA2X2 g91135(.A (n_2631), .B (n_2508), .Q (n_2710));
  NO2X2 g91137(.A (n_2623), .B (n_2277), .Q (n_2729));
  OR2X4 g91138(.A (n_2623), .B (n_2622), .Q (n_2728));
  OR2X2 g91140(.A (n_2623), .B (n_2593), .Q (n_2724));
  NO3X1 g91141(.A (n_2483), .B (store_type), .C (n_852), .Q (n_2721));
  INX1 g91143(.A (n_2690), .Q (n_2689));
  INX1 g91144(.A (n_2688), .Q (n_2687));
  NO2X2 g91145(.A (n_2633), .B (csr_mcause_code[3]), .Q
       (irq_software_response));
  AND2X1 g91146(.A (n_2632), .B (csr_mcause_code[3]), .Q
       (irq_external_response));
  NA2X2 g91147(.A (n_2621), .B (instruction[24]), .Q (n_2683));
  AND3X1 g91148(.A (n_2574), .B (n_2419), .C (csr_mcause_code[2]), .Q
       (irq_timer_response));
  NO2I1X1 g91149(.B (n_4451), .AN (n_8049), .Q (n_2709));
  NA2I1X1 g91150(.B (n_8035), .AN (n_4439), .Q (n_2708));
  AND2X1 g91151(.A (n_8029), .B (n_4434), .Q (n_2707));
  NA2I1X1 g91152(.B (n_8031), .AN (n_4436), .Q (n_2706));
  NA2X1 g91153(.A (n_8047), .B (n_4449), .Q (n_2705));
  NA2I1X1 g91154(.B (n_8041), .AN (n_4444), .Q (n_2704));
  AND2X1 g91155(.A (n_8040), .B (n_4443), .Q (n_2703));
  NA2X1 g91156(.A (n_8042), .B (n_4445), .Q (n_2702));
  NO2I1X1 g91157(.B (n_4450), .AN (n_8048), .Q (n_2701));
  NO2X4 g91158(.A (n_2621), .B (instruction[24]), .Q (n_8164));
  NA2X1 g91159(.A (n_8033), .B (n_4437), .Q (n_2700));
  AND2X1 g91160(.A (n_8046), .B (n_4448), .Q (n_2699));
  AND2X1 g91161(.A (n_8043), .B (n_4446), .Q (n_2698));
  NA2I1X1 g91162(.B (n_8037), .AN (n_4441), .Q (n_2697));
  NO2I1X1 g91163(.B (n_4442), .AN (n_8039), .Q (n_2696));
  NA2X1 g91164(.A (n_8034), .B (n_4438), .Q (n_2695));
  NA2X1 g91165(.A (n_8028), .B (n_4433), .Q (n_2694));
  NA2X1 g91166(.A (n_8030), .B (n_4435), .Q (n_2693));
  NA2I1X1 g91167(.B (n_8036), .AN (n_4440), .Q (n_2692));
  NA2X1 g91168(.A (n_8045), .B (n_4447), .Q (n_2691));
  NO2I1X1 g91169(.B (n_2630), .AN (csr_mcause_code[3]), .Q (n_2690));
  AND2X1 g91170(.A (n_2639), .B (csr_mcause_code[3]), .Q (n_2688));
  NO2X1 g91171(.A (n_2630), .B (csr_mcause_code[3]), .Q (n_2686));
  NO2I1X1 g91172(.B (csr_mcause_code[3]), .AN (n_2639), .Q (n_2685));
  NA2I1X4 g91173(.B (n_2613), .AN (n_2606), .Q (n_2684));
  AND2X1 g91174(.A (\rs1_data[21]_39616 ), .B (n_2589), .Q (n_2682));
  MU2IX1 g91176(.S (alu_sra_result[31]), .IN0 (n_8160), .IN1 (n_8161),
       .Q (n_2680));
  ON21X1 g91178(.A (\rs1_data[15]_39556 ), .B (n_2476), .C (n_2310), .Q
       (n_2678));
  NO2X1 g91180(.A (n_2528), .B (n_2590), .Q (n_2676));
  NO2X1 g91184(.A (n_2426), .B (n_2588), .Q (n_2672));
  NA2X1 g91185(.A (\rs1_data[30]_39526 ), .B (n_2589), .Q (n_2671));
  NA2X1 g91186(.A (alu_sra_result[31]), .B (n_2589), .Q (n_2670));
  NA2X1 g91187(.A (n_6135), .B (n_2589), .Q (n_2669));
  NA2X1 g91188(.A (\rs1_data[29]_39416 ), .B (n_2589), .Q (n_2668));
  NA2X1 g91189(.A (\rs1_data[22]_39626 ), .B (n_2589), .Q (n_2667));
  NA2X1 g91190(.A (\rs1_data[26]_39356 ), .B (n_2589), .Q (n_2666));
  NA2X1 g91192(.A (n_6136), .B (n_2589), .Q (n_2664));
  NA2X1 g91194(.A (\rs1_data[13]_39536 ), .B (n_2589), .Q (n_2662));
  AND2X1 g91196(.A (\rs1_data[19]_39596 ), .B (n_2589), .Q (n_2661));
  AN21X1 g91197(.A (n_501), .B (n_2477), .C (n_2590), .Q (n_2660));
  NA2X1 g91198(.A (\rs1_data[6]_39456 ), .B (n_2589), .Q (n_2659));
  NA2X1 g91199(.A (\rs1_data[7]_39466 ), .B (n_2589), .Q (n_2658));
  NA2X1 g91202(.A (\rs1_data[12]_39516 ), .B (n_2589), .Q (n_2656));
  ON21X1 g91203(.A (n_6132), .B (n_2476), .C (n_2310), .Q (n_2655));
  NA2X2 g91204(.A (n_6123), .B (n_2589), .Q (n_2654));
  NA2X2 g91205(.A (\rs1_data[4]_39436 ), .B (n_2589), .Q (n_2653));
  NA2X2 g91208(.A (n_8360), .B (n_2310), .Q (n_2651));
  NA2X1 g91209(.A (n_8366), .B (n_2589), .Q (n_2650));
  NA2X1 g91210(.A (n_2306), .B (n_2589), .Q (n_2649));
  NA2X1 g91211(.A (\rs1_data[9]_39486 ), .B (n_2589), .Q (n_2648));
  NA2X2 g91212(.A (n_2580), .B (n_2506), .Q (n_2647));
  AN21X1 g91213(.A (n_2437), .B (n_2506), .C (n_2310), .Q (n_2646));
  NA2X1 g91214(.A (n_2437), .B (n_2311), .Q (n_2645));
  NA2X1 g91215(.A (n_7681), .B (n_2311), .Q (n_2644));
  NO2X1 g91218(.A (n_2579), .B (n_2507), .Q (n_2642));
  AND2X1 g91219(.A (n_7692), .B (n_2311), .Q (n_2641));
  NA2X1 g91220(.A (n_2587), .B (n_7248), .Q (n_2640));
  INX1 g91221(.A (n_2637), .Q (n_2638));
  INX1 g91222(.A (n_2632), .Q (n_2633));
  INX1 g91223(.A (n_2627), .Q (n_2626));
  BUX2 g91225(.A (n_2621), .Q (n_2622));
  INX4 g91227(.A (n_2620), .Q (n_2619));
  INX2 g91238(.A (n_2314), .Q (n_2313));
  INX1 g91240(.A (n_2312), .Q (n_2615));
  BUX3 g91244(.A (n_2614), .Q (n_2312));
  NA2X1 g91246(.A (n_2601), .B (n_2424), .Q (n_2613));
  NA2X1 g91248(.A (n_2587), .B (n_6535), .Q (n_2611));
  NA2X1 g91250(.A (n_2597), .B (n_2595), .Q (n_2609));
  NO2X2 g91253(.A (n_2601), .B (n_2424), .Q (n_2606));
  NA2X1 g91255(.A (n_2309), .B (n_8053), .Q (n_2604));
  AND2X1 g91256(.A (n_2309), .B (n_8054), .Q (n_2603));
  NO2X1 g91257(.A (n_2573), .B (csr_mcause_code[2]), .Q (n_2639));
  NO2X1 g91259(.A (n_2593), .B (n_2513), .Q (n_2637));
  NO3X1 g91260(.A (n_2275), .B (n_2501), .C (n_2491), .Q (n_2636));
  AND2X1 g91261(.A (n_8162), .B (n_2571), .Q (n_2635));
  NA2X1 g91264(.A (n_2495), .B (n_2601), .Q (n_2634));
  NO2I1X1 g91268(.B (csr_mcause_code[2]), .AN (n_2574), .Q (n_2632));
  NO2X2 g91269(.A (n_2600), .B (n_2593), .Q (n_2631));
  NA2X1 g91270(.A (n_2572), .B (csr_mcause_code[2]), .Q (n_2630));
  ON311X1 g91273(.A (n_6082), .B (current_state[3]), .C (n_2465), .D
       (n_7249), .E (n_8078), .Q (n_2628));
  NA2X1 g91286(.A (n_8163), .B (n_2571), .Q (n_2627));
  NA2X4 g91287(.A (n_2591), .B (n_8570), .Q (n_2625));
  NA3I1X4 g91288(.B (n_8570), .C (n_8486), .AN (n_2264), .Q (n_2623));
  NA2X4 g91289(.A (n_2489), .B (n_2601), .Q (n_2621));
  NA2X4 g91291(.A (n_2598), .B (n_2591), .Q (n_2620));
  NA2X2 g91292(.A (n_2598), .B (n_2508), .Q (n_2314));
  INX1 g91293(.A (n_2504), .Q (n_2602));
  INX4 g91294(.A (n_2478), .Q (n_2601));
  INX1 g91298(.A (n_2593), .Q (n_2592));
  INX1 g91300(.A (n_2589), .Q (n_2588));
  INX2 g91301(.A (n_2587), .Q (n_2586));
  NO2X1 g91302(.A (n_7682), .B (n_2505), .Q (n_2585));
  NO2X2 g91304(.A (\rs1_data[3]_39426 ), .B (n_8309), .Q (n_2584));
  NO2X2 g91305(.A (\rs1_data[1]_39396 ), .B (n_8309), .Q (n_2583));
  NO2X1 g91306(.A (n_7680), .B (n_2505), .Q (n_2582));
  NO2X2 g91307(.A (n_6123), .B (n_8309), .Q (n_2581));
  NA2X2 g91308(.A (n_2438), .B (n_8158), .Q (n_2580));
  NO2X1 g91309(.A (n_7692), .B (n_2505), .Q (n_2579));
  AN21X1 g91310(.A (n_2483), .B (n_8163), .C (jal_type), .Q (n_2578));
  NO2I1X1 g91311(.B (n_8306), .AN (n_2518), .Q (n_2577));
  NO2X2 g91312(.A (\rs1_data[4]_39436 ), .B (n_8309), .Q (n_2576));
  NO2X2 g91313(.A (n_2516), .B (n_2512), .Q (n_2600));
  NO2X1 g91314(.A (n_2522), .B (n_2305), .Q (n_2599));
  NO2X4 g91315(.A (n_2517), .B (n_2277), .Q (n_2598));
  NA2I1X1 g91317(.B (n_8484), .AN (n_8160), .Q (n_2597));
  NA2I1X1 g91318(.B (store_type), .AN (n_2514), .Q (n_2596));
  NO3X1 g91319(.A (n_2275), .B (n_8359), .C (n_8482), .Q (n_2595));
  NA2X1 g91321(.A (n_2518), .B (n_2502), .Q (n_8073));
  NA2X2 g91322(.A (n_2521), .B (n_2305), .Q (n_2593));
  NO2X4 g91323(.A (n_2275), .B (instruction[24]), .Q (n_2591));
  OR2X4 g91324(.A (n_2507), .B (n_8158), .Q (n_2590));
  AND2X4 g91325(.A (n_2276), .B (n_2416), .Q (n_2589));
  NO2X4 g91326(.A (n_2277), .B (instruction[24]), .Q (n_2587));
  INX1 g91327(.A (n_2572), .Q (n_2573));
  INX1 g91328(.A (n_2571), .Q (n_2570));
  INX1 g91341(.A (n_8207), .Q (n_2309));
  AND2X1 g91343(.A (n_2503), .B (irq_fast[15]), .Q (n_2567));
  AND2X1 g91344(.A (n_2503), .B (irq_fast[3]), .Q (n_2566));
  AND2X1 g91345(.A (n_2503), .B (irq_fast[9]), .Q (n_2565));
  NA2X1 g91346(.A (n_8224), .B (n_2503), .Q (n_8167));
  AND2X1 g91347(.A (n_2503), .B (irq_fast[7]), .Q (n_2564));
  AND2X1 g91348(.A (n_2503), .B (irq_fast[5]), .Q (n_2563));
  AND2X1 g91349(.A (n_2503), .B (irq_fast[1]), .Q (n_2562));
  AND2X1 g91350(.A (n_2503), .B (irq_fast[4]), .Q (n_2561));
  AND2X1 g91351(.A (n_2503), .B (irq_fast[6]), .Q (n_2560));
  AND2X1 g91352(.A (n_2503), .B (irq_fast[2]), .Q (n_2559));
  AND2X1 g91353(.A (n_2503), .B (irq_fast[13]), .Q (n_2558));
  AND2X1 g91354(.A (n_2503), .B (irq_fast[0]), .Q (n_2557));
  AND2X1 g91355(.A (n_2503), .B (irq_timer), .Q (n_2556));
  AND2X1 g91356(.A (n_2503), .B (irq_fast[14]), .Q (n_2555));
  AND2X1 g91357(.A (n_2503), .B (irq_fast[11]), .Q (n_2554));
  AND2X1 g91358(.A (n_2503), .B (irq_fast[8]), .Q (n_2553));
  AND2X1 g91359(.A (n_2503), .B (irq_software), .Q (n_2552));
  AND2X1 g91360(.A (n_2503), .B (irq_external), .Q (n_2551));
  AND2X1 g91361(.A (n_2503), .B (irq_fast[10]), .Q (n_2550));
  AND2X1 g91362(.A (n_2503), .B (irq_fast[12]), .Q (n_2549));
  NO3X1 g91363(.A (n_2480), .B (csr_mcause_code[4]), .C (n_8078), .Q
       (n_2574));
  NO2I1X1 g91364(.B (n_8078), .AN (csr_mcause_code[4]), .Q (n_2572));
  NO2X1 g91365(.A (n_7714), .B (reset_internal_39074), .Q (n_2571));
  NO2X1 g91366(.A (n_2493), .B (n_8078), .Q (n_2569));
  NO2X1 g91367(.A (n_2492), .B (n_8078), .Q (n_2568));
  NA2X4 g91368(.A (n_7714), .B (n_2503), .Q (n_8207));
  NO2X1 g91370(.A (n_6149), .B (n_2476), .Q (n_2546));
  NO2X1 g91371(.A (n_6136), .B (n_2476), .Q (n_2545));
  NO2X1 g91372(.A (\rs1_data[26]_39356 ), .B (n_2476), .Q (n_2544));
  NO2X1 g91373(.A (alu_sra_result[31]), .B (n_2476), .Q (n_2543));
  NO2X1 g91374(.A (\rs1_data[23]_39326 ), .B (n_2476), .Q (n_2542));
  NO2X1 g91375(.A (n_6135), .B (n_2476), .Q (n_2541));
  NO2X1 g91376(.A (\rs1_data[22]_39626 ), .B (n_2476), .Q (n_2540));
  NO2X1 g91377(.A (\rs1_data[29]_39416 ), .B (n_2476), .Q (n_2539));
  NO2X1 g91378(.A (\rs1_data[30]_39526 ), .B (n_2476), .Q (n_2538));
  NO2X1 g91379(.A (\rs1_data[10]_39496 ), .B (n_2476), .Q (n_2537));
  NO2X1 g91380(.A (\rs1_data[11]_39506 ), .B (n_2476), .Q (n_2536));
  NO2X1 g91381(.A (\rs1_data[13]_39536 ), .B (n_2476), .Q (n_2535));
  NO2X1 g91382(.A (\rs1_data[24]_39336 ), .B (n_2476), .Q (n_2534));
  NO2X1 g91383(.A (\rs1_data[14]_39546 ), .B (n_2476), .Q (n_2533));
  NO2X1 g91384(.A (n_6141), .B (n_2476), .Q (n_2532));
  NO2X2 g91385(.A (\rs1_data[7]_39466 ), .B (n_2476), .Q (n_2531));
  NO2X1 g91386(.A (\rs1_data[21]_39616 ), .B (n_2476), .Q (n_2530));
  NO2X2 g91387(.A (\rs1_data[6]_39456 ), .B (n_2476), .Q (n_2529));
  NO2X1 g91388(.A (\rs1_data[19]_39596 ), .B (n_2476), .Q (n_2528));
  NO2X1 g91389(.A (\rs1_data[12]_39516 ), .B (n_2476), .Q (n_2527));
  NO2X1 g91390(.A (n_6127), .B (n_2476), .Q (n_2526));
  NO2X1 g91392(.A (\rs1_data[9]_39486 ), .B (n_2476), .Q (n_2524));
  NO2X1 g91393(.A (n_8366), .B (n_2476), .Q (n_2523));
  OR2X4 g91394(.A (n_2483), .B (jal_type), .Q (n_2548));
  INX1 g91396(.A (n_2521), .Q (n_2522));
  INX2 g91397(.A (n_2516), .Q (n_2517));
  INX1 g91398(.A (n_2515), .Q (n_8301));
  INX1 g91399(.A (n_2512), .Q (n_2513));
  INX1 g91400(.A (n_8159), .Q (n_2511));
  INX1 g91401(.A (n_2508), .Q (n_2509));
  INX1 g91402(.A (n_2507), .Q (n_2506));
  INX1 g91404(.A (n_2505), .Q (n_8158));
  INX1 g91405(.A (n_960), .Q (n_7249));
  INX1 g91406(.A (n_2503), .Q (reset_internal_39074));
  NO3X1 g91407(.A (n_2466), .B (instruction[3]), .C (instruction[2]),
       .Q (n_2502));
  NA3X1 g91408(.A (n_8484), .B (n_8482), .C (instruction[24]), .Q
       (n_2501));
  NA2I1X1 g91409(.B (branch_type), .AN (n_2308), .Q (n_2500));
  NA3I1X1 g91412(.B (system_type), .C (n_8163), .AN (n_8310), .Q
       (n_2520));
  NO3X1 g91415(.A (\instruction[5]_40251 ), .B (instruction[6]), .C
       (instruction[4]), .Q (n_2518));
  NO2X4 g91416(.A (n_8359), .B (n_2463), .Q (n_2516));
  NO2X1 g91417(.A (n_2481), .B (\instruction[14]_40189 ), .Q (n_2515));
  NA2X1 g91418(.A (n_2476), .B (n_2416), .Q (n_2514));
  NO2X4 g91419(.A (n_2467), .B (n_2491), .Q (n_2512));
  AND2X1 g91420(.A (n_7303), .B (n_2416), .Q (n_8162));
  NO2X1 g91423(.A (n_2481), .B (n_2416), .Q (n_8159));
  NA2X4 g91425(.A (n_2478), .B (n_2464), .Q (n_2510));
  NO4I1X4 g91426(.B (instruction[24]), .C (n_8486), .D (n_8485), .AN
       (n_8480), .Q (n_2508));
  NA2I1X2 g91427(.B (n_2481), .AN (n_7302), .Q (n_2507));
  NA2X2 g91428(.A (n_2308), .B (n_8676), .Q (n_8309));
  NA3I1X1 g91429(.B (n_2496), .C (n_6082), .AN (current_state[3]), .Q
       (n_8078));
  NA2X2 g91430(.A (n_2477), .B (\instruction[14]_40189 ), .Q (n_2505));
  AO21X1 g91431(.A (\instruction[8]_40127 ), .B (\instruction[7]_39642
       ), .C (n_2488), .Q (n_2504));
  NO2X2 g91433(.A (reset_reg), .B (reset), .Q (n_2503));
  INX1 g91435(.A (n_2492), .Q (n_2493));
  INX1 g91437(.A (n_2489), .Q (n_2490));
  INX1 g91438(.A (n_2480), .Q (n_2479));
  INCX12 g91441(.A (n_2477), .Q (n_2476));
  NA2X1 g91444(.A (n_7689), .B (n_2303), .Q (n_2472));
  NA2X2 g91456(.A (n_2421), .B (n_8482), .Q (n_2467));
  NA2X1 g91464(.A (instruction[0]), .B (instruction[1]), .Q (n_2466));
  NA2I1X0 g91465(.B (current_state[0]), .AN (current_state[1]), .Q
       (n_2465));
  NA2X1 g91466(.A (n_2431), .B (n_2415), .Q (n_2464));
  NO2X2 g91468(.A (n_8480), .B (n_8485), .Q (n_2498));
  NO2X1 g91469(.A (n_8302), .B (n_8303), .Q (n_2497));
  NO2X1 g91470(.A (current_state[0]), .B (current_state[1]), .Q
       (n_2496));
  NO2X1 g91471(.A (n_2424), .B (instruction[23]), .Q (n_2495));
  NA2X1 g91473(.A (n_8051), .B (csr_mcause_interrupt_flag), .Q
       (n_2492));
  NA2X2 g91474(.A (n_8484), .B (n_8482), .Q (n_2463));
  NA2X4 g91475(.A (instruction[28]), .B (n_8481), .Q (n_2491));
  NO2X4 g91476(.A (instruction[23]), .B (instruction[22]), .Q (n_2489));
  NO2X1 g91477(.A (\instruction[8]_40127 ), .B (\instruction[7]_39642
       ), .Q (n_2488));
  NO2X1 g91478(.A (n_4674), .B (n_8304), .Q (n_2487));
  NO2I1X1 g91479(.B (csr_mcause_code[1]), .AN (csr_mcause_code[0]), .Q
       (n_2486));
  NO2I1X1 g91480(.B (csr_mcause_code[0]), .AN (csr_mcause_code[1]), .Q
       (n_2485));
  NA2X1 g91481(.A (n_8157), .B (n_2390), .Q (n_2484));
  NO2X1 g91482(.A (n_8305), .B (n_8308), .Q (n_2483));
  NO2X1 g91483(.A (csr_mcause_code[0]), .B (csr_mcause_code[1]), .Q
       (n_2482));
  NA2I1X1 g91485(.B (n_8487), .AN (n_8676), .Q (n_2481));
  NA2X1 g91486(.A (csr_mcause_code[0]), .B (csr_mcause_code[1]), .Q
       (n_2480));
  NA2I1X4 g91488(.B (n_2414), .AN (instruction[21]), .Q (n_2478));
  NO2X1 g91489(.A (flush_37557), .B (n_7714), .Q (n_7882));
  AND2X2 g91490(.A (n_8487), .B (n_8676), .Q (n_2477));
  NO2X1 g91491(.A (n_7714), .B (reset), .Q (n_2475));
  NO2X1 g91492(.A (n_2390), .B (reset), .Q (n_2474));
  INX1 g91545(.A (n_7685), .Q (n_2462));
  INX1 g91546(.A (n_7242), .Q (n_2461));
  INX1 g91548(.A (n_7693), .Q (n_2460));
  INX1 g91549(.A (n_7670), .Q (n_2459));
  INX1 g91550(.A (n_8260), .Q (n_2458));
  INX1 g91551(.A (n_8257), .Q (n_2457));
  INX1 g91552(.A (n_6562), .Q (n_2456));
  INX1 g91553(.A (n_7215), .Q (n_2455));
  INX1 g91554(.A (n_6438), .Q (n_2454));
  INX1 g91555(.A (n_6436), .Q (n_2453));
  INX1 g91556(.A (n_6411), .Q (n_2452));
  INX1 g91557(.A (n_6905), .Q (n_2451));
  INX1 g91558(.A (n_6440), .Q (n_2450));
  INX1 g91559(.A (n_6409), .Q (n_2449));
  INX1 g91560(.A (n_6564), .Q (n_2448));
  INX1 g91561(.A (n_6362), .Q (n_2447));
  INX1 g91562(.A (n_6405), .Q (n_2446));
  INX1 g91563(.A (n_7217), .Q (n_2445));
  INX1 g91564(.A (n_6560), .Q (n_2444));
  INX1 g91565(.A (program_counter[2]), .Q (n_7925));
  INX1 g91567(.A (\instruction[11]_40312 ), .Q (n_2442));
  INX1 g91568(.A (\instruction[9]_40095 ), .Q (n_2441));
  INX1 g91569(.A (\instruction[10]_40063 ), .Q (n_2440));
  INX1 g91570(.A (n_7682), .Q (n_2439));
  INX2 g91571(.A (n_7681), .Q (n_2438));
  INX2 g91573(.A (\rs1_data[25]_39346 ), .Q (n_501));
  INX1 g91575(.A (\rs1_data[15]_39556 ), .Q (n_2435));
  INX3 g91580(.A (n_6121), .Q (n_2433));
  INX1 g91583(.A (\rs1_data[23]_39326 ), .Q (n_2432));
  BUX2 g91584(.A (instruction[21]), .Q (n_2431));
  INX2 g91588(.A (\rs1_data[11]_39506 ), .Q (n_2429));
  INX1 g91590(.A (\rs1_data[6]_39456 ), .Q (n_2428));
  INX2 g91592(.A (\rs1_data[10]_39496 ), .Q (n_2426));
  INX1 g91594(.A (\rs1_data[14]_39546 ), .Q (n_2425));
  INX2 g91595(.A (instruction[22]), .Q (n_2424));
  INX1 g91596(.A (n_6135), .Q (n_2423));
  INX2 g91601(.A (n_8484), .Q (n_2421));
  INX1 g91602(.A (alu_sra_result[31]), .Q (n_2420));
  INX1 g91604(.A (csr_mcause_code[3]), .Q (n_2419));
  INX1 g91605(.A (n_8163), .Q (n_2418));
  INX1 g91606(.A (\instruction[7]_39642 ), .Q (n_2417));
  INX1 g91607(.A (\instruction[14]_40189 ), .Q (n_2416));
  BUX2 g91613(.A (n_2415), .Q (n_2304));
  INX2 g91614(.A (n_2414), .Q (n_2415));
  INX4 g91615(.A (instruction[20]), .Q (n_2414));
  INX3 g91622(.A (n_2303), .Q (n_2258));
  INX3 g91643(.A (\instruction[5]_40251 ), .Q (n_2303));
  INX1 g91644(.A (n_6566), .Q (n_2411));
  INX1 g91645(.A (n_6407), .Q (n_2410));
  INX1 g91646(.A (n_6442), .Q (n_2409));
  INX1 g91647(.A (n_6903), .Q (n_2408));
  INX1 g91648(.A (n_6907), .Q (n_2407));
  INX1 g91649(.A (n_6901), .Q (n_2406));
  INX1 g91650(.A (n_6318), .Q (n_2405));
  INX1 g91651(.A (n_6312), .Q (n_2404));
  INX1 g91652(.A (n_6938), .Q (n_2403));
  INX1 g91653(.A (n_6936), .Q (n_2402));
  INX1 g91654(.A (n_6910), .Q (n_2401));
  INX1 g91655(.A (n_6911), .Q (n_2400));
  INX1 g91656(.A (n_6575), .Q (n_2399));
  INX1 g91657(.A (n_6574), .Q (n_2398));
  INX1 g91658(.A (n_6469), .Q (n_2397));
  INX1 g91659(.A (n_6451), .Q (n_2396));
  INX1 g91660(.A (n_6450), .Q (n_2395));
  INX1 g91661(.A (n_6467), .Q (n_2394));
  INX1 g91662(.A (n_6480), .Q (n_2393));
  INX1 g91663(.A (n_6483), .Q (n_2392));
  INX4 g91665(.A (flush_37557), .Q (n_7883));
  INX1 g91667(.A (n_7714), .Q (n_2390));
  INX1 fopt91668(.A (n_8566), .Q (n_957));
  INX6 fopt91681(.A (n_3151), .Q (n_2300));
  NA2X4 g52647(.A (n_1169), .B (n_3008), .Q (n_2298));
  OR2X4 g91683(.A (n_8526), .B (n_2682), .Q (n_7385));
  OR2X4 g91685(.A (n_3516), .B (n_2714), .Q (n_7633));
  NA3I1X1 g91686(.B (n_4385), .C (n_4379), .AN (n_2279), .Q (n_2297));
  NA2I1X2 g91687(.B (n_4316), .AN (n_2294), .Q (n_2296));
  OR2X2 g91688(.A (n_4279), .B (n_4204), .Q (n_2295));
  NA3I1X2 g91689(.B (n_4249), .C (n_4232), .AN (n_4278), .Q (n_2294));
  NA3I1X1 g91690(.B (n_8492), .C (n_2288), .AN (n_8493), .Q (n_2293));
  OR2X2 g91691(.A (n_4244), .B (n_4245), .Q (n_2292));
  NA2I1X1 g91693(.B (n_2268), .AN (n_4226), .Q (n_2290));
  MU2IX1 g91694(.S (n_8496), .IN0 (alu_operation_code_39112), .IN1
       (n_2326), .Q (n_8293));
  NA3I2X1 g91695(.C (n_4226), .AN (n_2380), .BN (n_2381), .Q (n_2289));
  NO3I1X1 g91696(.B (n_4201), .C (n_4174), .AN (n_4207), .Q (n_2288));
  NA2I1X1 g91698(.B (n_4238), .AN (n_4201), .Q (n_2286));
  NO3I1X1 g91699(.B (n_4227), .C (n_2378), .AN (n_4175), .Q (n_2285));
  NA2I1X1 g91700(.B (n_4204), .AN (n_2375), .Q (n_2284));
  MU2X2 g91701(.S (n_2258), .IN0 (n_7669), .IN1 (n_2368), .Q
       (alu_2nd_operand[22]));
  NA2I1X1 g91702(.B (\rs1_data[13]_39536 ), .AN (n_4132), .Q (n_2283));
  NO3I1X1 g91703(.B (\instruction[7]_39642 ), .C (n_3007), .AN
       (n_3179), .Q (n_2282));
  NA2I1X1 g91704(.B (n_2309), .AN (n_3182), .Q (n_8168));
  NA2I1X2 g91705(.B (n_2939), .AN (n_3005), .Q (n_2281));
  NA2I1X4 g91706(.B (n_3082), .AN (n_2857), .Q (n_2280));
  NO3I1X1 g91707(.B (n_2708), .C (n_4367), .AN (n_2695), .Q (n_2279));
  NA3I1X1 g91708(.B (n_3044), .C (n_2969), .AN (n_2316), .Q (n_2278));
  NO3I1X1 g91709(.B (n_8484), .C (n_2520), .AN (n_2595), .Q (n_7371));
  OR2X4 g91710(.A (n_2490), .B (n_2263), .Q (n_2277));
  NA2I1X1 g91711(.B (n_2481), .AN (n_7303), .Q (n_2276));
  NA2I1X2 g91712(.B (n_2498), .AN (n_8486), .Q (n_2275));
  NA2I1X2 g91713(.B (n_2368), .AN (\rs1_data[22]_39626 ), .Q (n_2274));
  NA2I1X1 g91714(.B (n_4127), .AN (\rs1_data[9]_39486 ), .Q (n_2273));
  NA2I1X2 g91715(.B (n_4118), .AN (\rs1_data[3]_39426 ), .Q (n_2272));
  NA2I1X1 g91716(.B (n_4124), .AN (n_6123), .Q (n_2271));
  NA2I1X1 g91718(.B (n_4152), .AN (\rs1_data[29]_39416 ), .Q (n_2269));
  NA2I1X1 g91719(.B (n_2363), .AN (\rs1_data[7]_39466 ), .Q (n_2268));
  NA2I1X1 g91720(.B (n_4151), .AN (\rs1_data[30]_39526 ), .Q (n_2267));
  NA2I1X1 g91721(.B (n_4150), .AN (n_6136), .Q (n_2266));
  NA2I1X1 g91722(.B (n_4132), .AN (\rs1_data[13]_39536 ), .Q (n_2265));
  NA2I1X2 g91723(.B (n_2498), .AN (instruction[24]), .Q (n_2264));
  NA2I1X2 g91724(.B (n_2415), .AN (n_2431), .Q (n_2263));
  NO3I2X1 g91726(.C (n_6082), .AN (n_2496), .BN (current_state[3]), .Q
       (n_960));
  INX2 g91730(.A (n_3060), .Q (n_2335));
  AND2X1 g91734(.A (n_3161), .B (n_7180), .Q (n_2343));
  AND2X1 g91736(.A (n_3382), .B (n_3504), .Q (n_2352));
  AND2X1 g91740(.A (n_3511), .B (n_3499), .Q (n_2347));
  AND2X1 g91746(.A (n_3700), .B (n_3701), .Q (n_2359));
  AND2X1 g91748(.A (n_3688), .B (n_3689), .Q (n_2360));
  AND2X1 g91750(.A (n_3440), .B (n_3380), .Q (n_2353));
  AND2X1 g91752(.A (n_3745), .B (n_3766), .Q (n_2361));
  AND6X1 g91754(.A (n_2870), .B (n_2872), .C (n_2998), .D (n_2933), .E
       (n_2835), .F (n_2776), .Q (n_2346));
  AND2X1 g91756(.A (n_3564), .B (n_3541), .Q (n_2357));
  INX2 g91768(.A (n_2856), .Q (n_2328));
  INX1 g91776(.A (n_7882), .Q (n_2307));
  NO2I1X1 g91786(.B (n_8487), .AN (n_8676), .Q (n_7303));
  OA21X1 g91788(.A (n_2537), .B (n_2590), .C (csr_data_out[10]), .Q
       (n_2345));
  INX2 g91790(.A (n_2272), .Q (n_2374));
  NO2I1X1 g91792(.B (n_4124), .AN (n_6123), .Q (n_2378));
  AND2X2 g91794(.A (n_2268), .B (n_4192), .Q (n_2383));
  INX1 g91796(.A (n_4170), .Q (n_2372));
  INX1 g91798(.A (n_4148), .Q (n_2371));
  INX1 g91800(.A (n_2369), .Q (n_2370));
  NO2I1X2 g91802(.B (n_2371), .AN (n_6149), .Q (n_2380));
  NO2I1X2 g91804(.B (n_2370), .AN (\rs1_data[21]_39616 ), .Q (n_2381));
  NO2I1X2 g91806(.B (n_4119), .AN (\rs1_data[1]_39396 ), .Q (n_2375));
  INX1 g91808(.A (n_4118), .Q (n_2365));
  NO2I1X1 g91810(.B (n_4127), .AN (\rs1_data[9]_39486 ), .Q (n_2377));
  NO2I1X2 g91812(.B (n_8619), .AN (\rs1_data[26]_39356 ), .Q (n_2379));
  INX2 g91814(.A (n_4119), .Q (n_2366));
  AND2X1 g91820(.A (n_2276), .B (\instruction[14]_40189 ), .Q (n_2311));
  INX2 g91822(.A (n_8659), .Q (n_2331));
  OR5X1 g91824(.A (n_2548), .B (n_4696), .C (n_2487), .D (n_2497), .E
       (n_852), .Q (n_2329));
  INX1 g91826(.A (n_2590), .Q (n_2310));
  NO2I1X2 g91828(.B (n_2367), .AN (\rs1_data[4]_39436 ), .Q (n_2373));
  NO2I1X1 g91830(.B (n_4251), .AN (n_4205), .Q (n_2287));
  AND2X2 g91832(.A (n_2269), .B (n_2266), .Q (n_2384));
  OA21X1 g91834(.A (n_4376), .B (n_2570), .C (n_2604), .Q (n_2389));
  INX2 g91836(.A (n_4382), .Q (n_2388));
  NA2I1X4 g91837(.B (n_2599), .AN (n_2623), .Q (n_2260));
  NA2I1X4 g91838(.B (n_2433), .AN (n_8309), .Q (n_2259));
  AND2X1 g91842(.A (n_3405), .B (n_3506), .Q (n_2351));
  AND2X1 g91844(.A (n_3450), .B (n_3424), .Q (n_2349));
  AND2X1 g91846(.A (n_3423), .B (n_3363), .Q (n_2348));
  OA21X1 g91848(.A (n_2514), .B (n_2515), .C (n_2571), .Q (n_2316));
  AND2X1 g91850(.A (n_6149), .B (n_2589), .Q (n_2320));
  AND2X1 g91852(.A (n_6141), .B (n_2589), .Q (n_2319));
  AND2X1 g91854(.A (n_6127), .B (n_2589), .Q (n_2318));
  NO2I1X2 g91856(.B (n_2372), .AN (\rs1_data[13]_39536 ), .Q (n_2382));
  AND2X1 g91858(.A (n_7303), .B (\instruction[14]_40189 ), .Q (n_8160));
  AND2X1 g91860(.A (n_2416), .B (n_8487), .Q (n_2308));
  NA3X1 g28110(.A (n_2237), .B (n_2242), .C (n_2253), .Q (n_2257));
  NA2X1 g28112(.A (n_2255), .B (n_2237), .Q (n_2256));
  NO2X1 g28114(.A (n_2235), .B (n_8216), .Q (n_2255));
  NO2X1 g28115(.A (n_2251), .B (n_8214), .Q (n_2254));
  NO3X1 g28116(.A (n_8209), .B (n_2238), .C (n_2250), .Q (n_2253));
  NA3X1 g28118(.A (n_2237), .B (n_2249), .C (n_2241), .Q (n_2252));
  OR6X1 g28120(.A (n_8215), .B (n_8222), .C (n_8221), .D (n_8223), .E
       (n_8365), .F (n_8219), .Q (n_2251));
  NA3I1X1 g28121(.B (n_2246), .C (n_18079_BAR), .AN (n_8218), .Q
       (n_2250));
  NO3X1 g28122(.A (n_8209), .B (n_8215), .C (n_2245), .Q (n_2249));
  OR3X1 g28123(.A (n_8219), .B (n_8218), .C (n_2244), .Q (n_2248));
  AN211X1 g28125(.A (n_7861), .B (n_7882), .C (n_2244), .D (n_8223), .Q
       (n_2246));
  NA2X1 g28126(.A (n_18082_BAR), .B (n_2239), .Q (n_2245));
  AND2X1 g28127(.A (take_trap_39229), .B (n_2240), .Q (n_2243));
  NO3I1X1 g28128(.B (n_8300), .C (n_2236), .AN (n_7371), .Q (n_2244));
  NO3X1 g28129(.A (n_8216), .B (n_8211), .C (n_8210), .Q (n_2242));
  NO3X1 g28130(.A (n_2238), .B (n_8213), .C (n_8222), .Q (n_2241));
  NO3I1X1 g28131(.B (n_7862), .C (n_7860), .AN (n_7882), .Q (n_2240));
  ON21X1 g28132(.A (n_7860), .B (n_7859), .C (n_7882), .Q (n_2239));
  OR2X1 g28133(.A (n_8221), .B (n_8220), .Q (n_2238));
  NO2X1 g28134(.A (n_8214), .B (n_8212), .Q (n_2237));
  NA2X1 g28135(.A (n_8164), .B (n_7882), .Q (n_2236));
  OR5X1 g28138(.A (n_8211), .B (n_8215), .C (n_2248), .D (n_8213), .E
       (n_8217), .Q (n_2235));
  DFRQX1 \csr_mcause_reg[0] (.C (rc_gclk_199882), .D (n_2234), .Q
       (csr_mcause[0]));
  DFRQX1 \csr_mcause_reg[10] (.C (rc_gclk_199882), .D (n_147), .Q
       (csr_mcause[10]));
  DFRQX1 \csr_mcause_reg[11] (.C (rc_gclk_199882), .D (n_146), .Q
       (csr_mcause[11]));
  DFRQX1 \csr_mcause_reg[12] (.C (rc_gclk_199882), .D (n_145), .Q
       (csr_mcause[12]));
  DFRQX1 \csr_mcause_reg[13] (.C (rc_gclk_199882), .D (n_144), .Q
       (csr_mcause[13]));
  DFRQX1 \csr_mcause_reg[14] (.C (rc_gclk_199882), .D (n_143), .Q
       (csr_mcause[14]));
  DFRQX1 \csr_mcause_reg[15] (.C (rc_gclk_199882), .D (n_142), .Q
       (csr_mcause[15]));
  DFRQX1 \csr_mcause_reg[16] (.C (rc_gclk_199882), .D (n_141), .Q
       (csr_mcause[16]));
  DFRQX1 \csr_mcause_reg[17] (.C (rc_gclk_199882), .D (n_140), .Q
       (csr_mcause[17]));
  DFRQX1 \csr_mcause_reg[18] (.C (rc_gclk_199882), .D (n_139), .Q
       (csr_mcause[18]));
  DFRQX1 \csr_mcause_reg[19] (.C (rc_gclk_199882), .D (n_138), .Q
       (csr_mcause[19]));
  DFRQX1 \csr_mcause_reg[1] (.C (rc_gclk_199882), .D (n_2233), .Q
       (csr_mcause[1]));
  DFRQX1 \csr_mcause_reg[20] (.C (rc_gclk_199882), .D (n_137), .Q
       (csr_mcause[20]));
  DFRQX1 \csr_mcause_reg[21] (.C (rc_gclk_199882), .D (n_136), .Q
       (csr_mcause[21]));
  DFRQX1 \csr_mcause_reg[22] (.C (rc_gclk_199882), .D (n_135), .Q
       (csr_mcause[22]));
  DFRQX1 \csr_mcause_reg[23] (.C (rc_gclk_199882), .D (n_134), .Q
       (csr_mcause[23]));
  DFRQX1 \csr_mcause_reg[24] (.C (rc_gclk_199882), .D (n_133), .Q
       (csr_mcause[24]));
  DFRQX1 \csr_mcause_reg[25] (.C (rc_gclk_199882), .D (n_132), .Q
       (csr_mcause[25]));
  DFRQX1 \csr_mcause_reg[26] (.C (rc_gclk_199882), .D (n_131), .Q
       (csr_mcause[26]));
  DFRQX1 \csr_mcause_reg[27] (.C (rc_gclk_199882), .D (n_130), .Q
       (csr_mcause[27]));
  DFRQX1 \csr_mcause_reg[28] (.C (rc_gclk_199882), .D (n_129), .Q
       (csr_mcause[28]));
  DFRQX1 \csr_mcause_reg[29] (.C (rc_gclk_199882), .D (n_128), .Q
       (csr_mcause[29]));
  DFRQX1 \csr_mcause_reg[2] (.C (rc_gclk_199882), .D (n_2232), .Q
       (csr_mcause[2]));
  DFRQX1 \csr_mcause_reg[30] (.C (rc_gclk_199882), .D (n_2231), .Q
       (csr_mcause[30]));
  DFRQX1 \csr_mcause_reg[31] (.C (rc_gclk_199882), .D (n_2230), .Q
       (csr_mcause[31]));
  DFRQX1 \csr_mcause_reg[3] (.C (rc_gclk_199882), .D (n_2229), .Q
       (csr_mcause[3]));
  DFRQX1 \csr_mcause_reg[4] (.C (rc_gclk_199882), .D (n_2228), .Q
       (csr_mcause[4]));
  DFRQX1 \csr_mcause_reg[5] (.C (rc_gclk_199882), .D (n_127), .Q
       (csr_mcause[5]));
  DFRQX1 \csr_mcause_reg[6] (.C (rc_gclk_199882), .D (n_126), .Q
       (csr_mcause[6]));
  DFRQX1 \csr_mcause_reg[7] (.C (rc_gclk_199882), .D (n_114), .Q
       (csr_mcause[7]));
  DFRQX1 \csr_mcause_reg[8] (.C (rc_gclk_199882), .D (n_125), .Q
       (csr_mcause[8]));
  DFRQX1 \csr_mcause_reg[9] (.C (rc_gclk_199882), .D (n_124), .Q
       (csr_mcause[9]));
  DFRQX1 \csr_mscratch_reg[0] (.C (rc_gclk_199966), .D (n_2063), .Q
       (csr_mscratch[0]));
  DFRQX1 \csr_mscratch_reg[10] (.C (rc_gclk_199966), .D (n_147), .Q
       (csr_mscratch[10]));
  DFRQX1 \csr_mscratch_reg[11] (.C (rc_gclk_199966), .D (n_146), .Q
       (csr_mscratch[11]));
  DFRQX1 \csr_mscratch_reg[12] (.C (rc_gclk_199966), .D (n_145), .Q
       (csr_mscratch[12]));
  DFRQX1 \csr_mscratch_reg[13] (.C (rc_gclk_199966), .D (n_144), .Q
       (csr_mscratch[13]));
  DFRQX1 \csr_mscratch_reg[14] (.C (rc_gclk_199966), .D (n_143), .Q
       (csr_mscratch[14]));
  DFRQX1 \csr_mscratch_reg[15] (.C (rc_gclk_199966), .D (n_142), .Q
       (csr_mscratch[15]));
  DFRQX1 \csr_mscratch_reg[16] (.C (rc_gclk_199966), .D (n_141), .Q
       (csr_mscratch[16]));
  DFRQX1 \csr_mscratch_reg[17] (.C (rc_gclk_199966), .D (n_140), .Q
       (csr_mscratch[17]));
  DFRQX1 \csr_mscratch_reg[18] (.C (rc_gclk_199966), .D (n_139), .Q
       (csr_mscratch[18]));
  DFRQX1 \csr_mscratch_reg[19] (.C (rc_gclk_199966), .D (n_138), .Q
       (csr_mscratch[19]));
  DFRQX1 \csr_mscratch_reg[1] (.C (rc_gclk_199966), .D (n_2062), .Q
       (csr_mscratch[1]));
  DFRQX1 \csr_mscratch_reg[20] (.C (rc_gclk_199966), .D (n_137), .Q
       (csr_mscratch[20]));
  DFRQX1 \csr_mscratch_reg[21] (.C (rc_gclk_199966), .D (n_136), .Q
       (csr_mscratch[21]));
  DFRQX1 \csr_mscratch_reg[22] (.C (rc_gclk_199966), .D (n_135), .Q
       (csr_mscratch[22]));
  DFRQX1 \csr_mscratch_reg[23] (.C (rc_gclk_199966), .D (n_134), .Q
       (csr_mscratch[23]));
  DFRQX1 \csr_mscratch_reg[24] (.C (rc_gclk_199966), .D (n_133), .Q
       (csr_mscratch[24]));
  DFRQX1 \csr_mscratch_reg[25] (.C (rc_gclk_199966), .D (n_132), .Q
       (csr_mscratch[25]));
  DFRQX1 \csr_mscratch_reg[26] (.C (rc_gclk_199966), .D (n_131), .Q
       (csr_mscratch[26]));
  DFRQX1 \csr_mscratch_reg[27] (.C (rc_gclk_199966), .D (n_130), .Q
       (csr_mscratch[27]));
  DFRQX1 \csr_mscratch_reg[28] (.C (rc_gclk_199966), .D (n_129), .Q
       (csr_mscratch[28]));
  DFRQX1 \csr_mscratch_reg[29] (.C (rc_gclk_199966), .D (n_128), .Q
       (csr_mscratch[29]));
  DFRQX1 \csr_mscratch_reg[2] (.C (rc_gclk_199966), .D (n_2061), .Q
       (csr_mscratch[2]));
  DFRQX1 \csr_mscratch_reg[30] (.C (rc_gclk_199966), .D (n_123), .Q
       (csr_mscratch[30]));
  DFRQX1 \csr_mscratch_reg[31] (.C (rc_gclk_199966), .D (n_2060), .Q
       (csr_mscratch[31]));
  DFRQX1 \csr_mscratch_reg[3] (.C (rc_gclk_199966), .D (n_2059), .Q
       (csr_mscratch[3]));
  DFRQX1 \csr_mscratch_reg[4] (.C (rc_gclk_199966), .D (n_2058), .Q
       (csr_mscratch[4]));
  DFRQX1 \csr_mscratch_reg[5] (.C (rc_gclk_199966), .D (n_127), .Q
       (csr_mscratch[5]));
  DFRQX1 \csr_mscratch_reg[6] (.C (rc_gclk_199966), .D (n_126), .Q
       (csr_mscratch[6]));
  DFRQX1 \csr_mscratch_reg[7] (.C (rc_gclk_199966), .D (n_114), .Q
       (csr_mscratch[7]));
  DFRQX1 \csr_mscratch_reg[8] (.C (rc_gclk_199966), .D (n_125), .Q
       (csr_mscratch[8]));
  DFRQX1 \csr_mscratch_reg[9] (.C (rc_gclk_199966), .D (n_124), .Q
       (csr_mscratch[9]));
  DFRQX1 \csr_mtval_reg[0] (.C (rc_gclk_199885), .D (n_2055), .Q
       (csr_mtval[0]));
  DFRQX1 \csr_mtval_reg[10] (.C (rc_gclk_199885), .D (n_2054), .Q
       (csr_mtval[10]));
  DFRQX1 \csr_mtval_reg[11] (.C (rc_gclk_199885), .D (n_2053), .Q
       (csr_mtval[11]));
  DFRQX1 \csr_mtval_reg[12] (.C (rc_gclk_199885), .D (n_2052), .Q
       (csr_mtval[12]));
  DFRQX1 \csr_mtval_reg[13] (.C (rc_gclk_199885), .D (n_2051), .Q
       (csr_mtval[13]));
  DFRQX1 \csr_mtval_reg[14] (.C (rc_gclk_199885), .D (n_2050), .Q
       (csr_mtval[14]));
  DFRQX1 \csr_mtval_reg[15] (.C (rc_gclk_199885), .D (n_2049), .Q
       (csr_mtval[15]));
  DFRQX1 \csr_mtval_reg[16] (.C (rc_gclk_199885), .D (n_2048), .Q
       (csr_mtval[16]));
  DFRQX1 \csr_mtval_reg[17] (.C (rc_gclk_199885), .D (n_2047), .Q
       (csr_mtval[17]));
  DFRQX1 \csr_mtval_reg[18] (.C (rc_gclk_199885), .D (n_2046), .Q
       (csr_mtval[18]));
  DFRQX1 \csr_mtval_reg[19] (.C (rc_gclk_199885), .D (n_2045), .Q
       (csr_mtval[19]));
  DFRQX1 \csr_mtval_reg[1] (.C (rc_gclk_199885), .D (n_2044), .Q
       (csr_mtval[1]));
  DFRQX1 \csr_mtval_reg[20] (.C (rc_gclk_199885), .D (n_2043), .Q
       (csr_mtval[20]));
  DFRQX1 \csr_mtval_reg[21] (.C (rc_gclk_199885), .D (n_2042), .Q
       (csr_mtval[21]));
  DFRQX1 \csr_mtval_reg[22] (.C (rc_gclk_199885), .D (n_2041), .Q
       (csr_mtval[22]));
  DFRQX1 \csr_mtval_reg[23] (.C (rc_gclk_199885), .D (n_2040), .Q
       (csr_mtval[23]));
  DFRQX1 \csr_mtval_reg[24] (.C (rc_gclk_199885), .D (n_2039), .Q
       (csr_mtval[24]));
  DFRQX1 \csr_mtval_reg[25] (.C (rc_gclk_199885), .D (n_2038), .Q
       (csr_mtval[25]));
  DFRQX1 \csr_mtval_reg[26] (.C (rc_gclk_199885), .D (n_2037), .Q
       (csr_mtval[26]));
  DFRQX1 \csr_mtval_reg[27] (.C (rc_gclk_199885), .D (n_2036), .Q
       (csr_mtval[27]));
  DFRQX1 \csr_mtval_reg[28] (.C (rc_gclk_199885), .D (n_2035), .Q
       (csr_mtval[28]));
  DFRQX1 \csr_mtval_reg[29] (.C (rc_gclk_199885), .D (n_2034), .Q
       (csr_mtval[29]));
  DFRQX1 \csr_mtval_reg[2] (.C (rc_gclk_199885), .D (n_2033), .Q
       (csr_mtval[2]));
  DFRQX1 \csr_mtval_reg[30] (.C (rc_gclk_199885), .D (n_2032), .Q
       (csr_mtval[30]));
  DFRQX1 \csr_mtval_reg[31] (.C (rc_gclk_199885), .D (n_2031), .Q
       (csr_mtval[31]));
  DFRQX1 \csr_mtval_reg[3] (.C (rc_gclk_199885), .D (n_2030), .Q
       (csr_mtval[3]));
  DFRQX1 \csr_mtval_reg[4] (.C (rc_gclk_199885), .D (n_2029), .Q
       (csr_mtval[4]));
  DFRQX1 \csr_mtval_reg[5] (.C (rc_gclk_199885), .D (n_2028), .Q
       (csr_mtval[5]));
  DFRQX1 \csr_mtval_reg[6] (.C (rc_gclk_199885), .D (n_2027), .Q
       (csr_mtval[6]));
  DFRQX1 \csr_mtval_reg[7] (.C (rc_gclk_199885), .D (n_2026), .Q
       (csr_mtval[7]));
  DFRQX1 \csr_mtval_reg[8] (.C (rc_gclk_199885), .D (n_2025), .Q
       (csr_mtval[8]));
  DFRQX1 \csr_mtval_reg[9] (.C (rc_gclk_199885), .D (n_2024), .Q
       (csr_mtval[9]));
  DFRQX4 \current_state_reg[0] (.C (rc_gclk_199995), .D (n_179), .Q
       (current_state[0]));
  DFRQX4 \current_state_reg[1] (.C (rc_gclk_199995), .D (n_2013), .Q
       (current_state[1]));
  DFRQX4 \current_state_reg[2] (.C (rc_gclk_199995), .D (n_2012), .Q
       (current_state[2]));
  DFRQX4 \current_state_reg[3] (.C (rc_gclk_199995), .D (n_2011), .Q
       (current_state[3]));
  DFRQX1 \prev_instruction_address_reg[0] (.C (rc_gclk), .D (n_1587),
       .Q (prev_instruction_address[0]));
  DFRQX1 \prev_instruction_reg[11] (.C (rc_gclk_199999), .D (n_1584),
       .Q (prev_instruction[11]));
  DFRQX4 prev_read_request_reg(.C (rc_gclk), .D (n_1553), .Q (n_8053));
  DFRQX1 \prev_rw_address_reg[0] (.C (rc_gclk), .D (n_184), .Q
       (prev_rw_address[0]));
  DFRQX1 \prev_rw_address_reg[10] (.C (rc_gclk), .D (n_1552), .Q
       (prev_rw_address[10]));
  DFRQX1 \prev_rw_address_reg[11] (.C (rc_gclk), .D (n_1551), .Q
       (prev_rw_address[11]));
  DFRQX1 \prev_rw_address_reg[12] (.C (rc_gclk), .D (n_1550), .Q
       (prev_rw_address[12]));
  DFRQX1 \prev_rw_address_reg[13] (.C (rc_gclk), .D (n_1549), .Q
       (prev_rw_address[13]));
  DFRQX1 \prev_rw_address_reg[14] (.C (rc_gclk), .D (n_1548), .Q
       (prev_rw_address[14]));
  DFRQX1 \prev_rw_address_reg[15] (.C (rc_gclk), .D (n_1547), .Q
       (prev_rw_address[15]));
  DFRQX1 \prev_rw_address_reg[16] (.C (rc_gclk), .D (n_1546), .Q
       (prev_rw_address[16]));
  DFRQX1 \prev_rw_address_reg[17] (.C (rc_gclk), .D (n_1545), .Q
       (prev_rw_address[17]));
  DFRQX1 \prev_rw_address_reg[18] (.C (rc_gclk), .D (n_1544), .Q
       (prev_rw_address[18]));
  DFRQX1 \prev_rw_address_reg[19] (.C (rc_gclk), .D (n_1543), .Q
       (prev_rw_address[19]));
  DFRQX1 \prev_rw_address_reg[1] (.C (rc_gclk), .D (n_183), .Q
       (prev_rw_address[1]));
  DFRQX1 \prev_rw_address_reg[20] (.C (rc_gclk), .D (n_1542), .Q
       (prev_rw_address[20]));
  DFRQX1 \prev_rw_address_reg[21] (.C (rc_gclk), .D (n_1541), .Q
       (prev_rw_address[21]));
  DFRQX1 \prev_rw_address_reg[22] (.C (rc_gclk), .D (n_1540), .Q
       (prev_rw_address[22]));
  DFRQX1 \prev_rw_address_reg[23] (.C (rc_gclk), .D (n_1539), .Q
       (prev_rw_address[23]));
  DFRQX1 \prev_rw_address_reg[24] (.C (rc_gclk), .D (n_1538), .Q
       (prev_rw_address[24]));
  DFRQX1 \prev_rw_address_reg[25] (.C (rc_gclk), .D (n_1537), .Q
       (prev_rw_address[25]));
  DFRQX1 \prev_rw_address_reg[26] (.C (rc_gclk), .D (n_1536), .Q
       (prev_rw_address[26]));
  DFRQX1 \prev_rw_address_reg[27] (.C (rc_gclk), .D (n_1535), .Q
       (prev_rw_address[27]));
  DFRQX1 \prev_rw_address_reg[28] (.C (rc_gclk), .D (n_1534), .Q
       (prev_rw_address[28]));
  DFRQX1 \prev_rw_address_reg[29] (.C (rc_gclk), .D (n_1533), .Q
       (prev_rw_address[29]));
  DFRQX1 \prev_rw_address_reg[2] (.C (rc_gclk), .D (n_1532), .Q
       (prev_rw_address[2]));
  DFRQX1 \prev_rw_address_reg[30] (.C (rc_gclk), .D (n_1531), .Q
       (prev_rw_address[30]));
  DFRQX1 \prev_rw_address_reg[31] (.C (rc_gclk), .D (n_1530), .Q
       (prev_rw_address[31]));
  DFRQX1 \prev_rw_address_reg[3] (.C (rc_gclk), .D (n_1529), .Q
       (prev_rw_address[3]));
  DFRQX1 \prev_rw_address_reg[4] (.C (rc_gclk), .D (n_1528), .Q
       (prev_rw_address[4]));
  DFRQX1 \prev_rw_address_reg[5] (.C (rc_gclk), .D (n_1527), .Q
       (prev_rw_address[5]));
  DFRQX1 \prev_rw_address_reg[6] (.C (rc_gclk), .D (n_1526), .Q
       (prev_rw_address[6]));
  DFRQX1 \prev_rw_address_reg[7] (.C (rc_gclk), .D (n_1525), .Q
       (prev_rw_address[7]));
  DFRQX1 \prev_rw_address_reg[8] (.C (rc_gclk), .D (n_1524), .Q
       (prev_rw_address[8]));
  DFRQX1 \prev_rw_address_reg[9] (.C (rc_gclk), .D (n_1523), .Q
       (prev_rw_address[9]));
  DFRQX1 \prev_write_data_reg[0] (.C (rc_gclk), .D (n_1522), .Q
       (prev_write_data[0]));
  DFRQX1 \prev_write_data_reg[10] (.C (rc_gclk), .D (n_1521), .Q
       (prev_write_data[10]));
  DFRQX1 \prev_write_data_reg[11] (.C (rc_gclk), .D (n_1520), .Q
       (prev_write_data[11]));
  DFRQX1 \prev_write_data_reg[12] (.C (rc_gclk), .D (n_1519), .Q
       (prev_write_data[12]));
  DFRQX1 \prev_write_data_reg[13] (.C (rc_gclk), .D (n_1518), .Q
       (prev_write_data[13]));
  DFRQX1 \prev_write_data_reg[14] (.C (rc_gclk), .D (n_1517), .Q
       (prev_write_data[14]));
  DFRQX1 \prev_write_data_reg[15] (.C (rc_gclk), .D (n_1516), .Q
       (prev_write_data[15]));
  DFRQX1 \prev_write_data_reg[16] (.C (rc_gclk), .D (n_1515), .Q
       (prev_write_data[16]));
  DFRQX1 \prev_write_data_reg[17] (.C (rc_gclk), .D (n_1514), .Q
       (prev_write_data[17]));
  DFRQX1 \prev_write_data_reg[18] (.C (rc_gclk), .D (n_1513), .Q
       (prev_write_data[18]));
  DFRQX1 \prev_write_data_reg[19] (.C (rc_gclk), .D (n_1512), .Q
       (prev_write_data[19]));
  DFRQX1 \prev_write_data_reg[1] (.C (rc_gclk), .D (n_1511), .Q
       (prev_write_data[1]));
  DFRQX1 \prev_write_data_reg[20] (.C (rc_gclk), .D (n_1510), .Q
       (prev_write_data[20]));
  DFRQX1 \prev_write_data_reg[21] (.C (rc_gclk), .D (n_1509), .Q
       (prev_write_data[21]));
  DFRQX1 \prev_write_data_reg[22] (.C (rc_gclk), .D (n_1508), .Q
       (prev_write_data[22]));
  DFRQX1 \prev_write_data_reg[23] (.C (rc_gclk), .D (n_1507), .Q
       (prev_write_data[23]));
  DFRQX1 \prev_write_data_reg[24] (.C (rc_gclk), .D (n_1506), .Q
       (prev_write_data[24]));
  DFRQX1 \prev_write_data_reg[25] (.C (rc_gclk), .D (n_1505), .Q
       (prev_write_data[25]));
  DFRQX1 \prev_write_data_reg[26] (.C (rc_gclk), .D (n_1504), .Q
       (prev_write_data[26]));
  DFRQX1 \prev_write_data_reg[27] (.C (rc_gclk), .D (n_1503), .Q
       (prev_write_data[27]));
  DFRQX1 \prev_write_data_reg[28] (.C (rc_gclk), .D (n_1502), .Q
       (prev_write_data[28]));
  DFRQX1 \prev_write_data_reg[29] (.C (rc_gclk), .D (n_1501), .Q
       (prev_write_data[29]));
  DFRQX1 \prev_write_data_reg[2] (.C (rc_gclk), .D (n_1500), .Q
       (prev_write_data[2]));
  DFRQX1 \prev_write_data_reg[30] (.C (rc_gclk), .D (n_1499), .Q
       (prev_write_data[30]));
  DFRQX1 \prev_write_data_reg[31] (.C (rc_gclk), .D (n_1498), .Q
       (prev_write_data[31]));
  DFRQX1 \prev_write_data_reg[3] (.C (rc_gclk), .D (n_1497), .Q
       (prev_write_data[3]));
  DFRQX1 \prev_write_data_reg[4] (.C (rc_gclk), .D (n_1496), .Q
       (prev_write_data[4]));
  DFRQX1 \prev_write_data_reg[5] (.C (rc_gclk), .D (n_1495), .Q
       (prev_write_data[5]));
  DFRQX1 \prev_write_data_reg[6] (.C (rc_gclk), .D (n_1494), .Q
       (prev_write_data[6]));
  DFRQX1 \prev_write_data_reg[7] (.C (rc_gclk), .D (n_1493), .Q
       (prev_write_data[7]));
  DFRQX1 \prev_write_data_reg[8] (.C (rc_gclk), .D (n_1492), .Q
       (prev_write_data[8]));
  DFRQX1 \prev_write_data_reg[9] (.C (rc_gclk), .D (n_1491), .Q
       (prev_write_data[9]));
  DFRQX1 \prev_write_strobe_reg[0] (.C (rc_gclk), .D (n_182), .Q
       (prev_write_strobe[0]));
  DFRQX1 \prev_write_strobe_reg[1] (.C (rc_gclk), .D (n_1489), .Q
       (prev_write_strobe[1]));
  DFRQX1 \prev_write_strobe_reg[2] (.C (rc_gclk), .D (n_1488), .Q
       (prev_write_strobe[2]));
  DFRQX1 \prev_write_strobe_reg[3] (.C (rc_gclk), .D (n_1487), .Q
       (prev_write_strobe[3]));
  NO2X1 g91861(.A (n_1453), .B (n_1), .Q (n_2234));
  NO2X1 g91862(.A (n_1452), .B (n_1), .Q (n_2233));
  NO2X1 g91863(.A (n_1451), .B (n_1), .Q (n_2232));
  AND2X1 g91864(.A (n_7376), .B (n_181), .Q (n_2231));
  NO2X1 g91865(.A (n_1450), .B (n_1), .Q (n_2230));
  NO2X1 g91866(.A (n_1449), .B (n_1), .Q (n_2229));
  NO2X1 g91867(.A (n_1448), .B (n_1), .Q (n_2228));
  AND2X1 g50215(.A (n_1446), .B (n_181), .Q (n_2227));
  NO2X1 g50154(.A (n_1445), .B (n_179), .Q (n_2226));
  NO2X1 g50149(.A (n_1444), .B (n_180), .Q (n_2225));
  NO2X1 g50158(.A (n_1443), .B (n_179), .Q (n_2224));
  NO2X1 g50153(.A (n_1442), .B (n_180), .Q (n_2223));
  NO2X1 g50150(.A (n_1441), .B (n_179), .Q (n_2222));
  NO2X1 g50144(.A (n_1440), .B (n_180), .Q (n_2221));
  NO2X1 g50199(.A (n_1439), .B (n_179), .Q (n_2220));
  NO2X1 g50140(.A (n_1438), .B (n_179), .Q (n_2219));
  NO2X1 g50133(.A (n_1437), .B (n_179), .Q (n_2218));
  NO2X1 g50127(.A (n_1436), .B (n_1), .Q (n_2217));
  NO2X1 g50197(.A (n_1435), .B (n_1), .Q (n_2216));
  NO2X1 g50141(.A (n_1434), .B (n_179), .Q (n_2215));
  NO2X1 g50134(.A (n_1433), .B (n_179), .Q (n_2214));
  NO2X1 g50126(.A (n_1432), .B (n_179), .Q (n_2213));
  NO2X1 g50122(.A (n_1431), .B (n_179), .Q (n_2212));
  NO2X1 g50135(.A (n_1430), .B (n_179), .Q (n_2211));
  NO2X1 g50128(.A (n_1429), .B (n_180), .Q (n_2210));
  NO2X1 g50123(.A (n_1428), .B (n_179), .Q (n_2209));
  NO2X1 g50118(.A (n_1427), .B (n_1), .Q (n_2208));
  NO2X1 g50119(.A (n_1426), .B (n_1), .Q (n_2207));
  NO2X1 g50116(.A (n_1425), .B (n_1), .Q (n_2206));
  NO2X1 g50195(.A (n_1424), .B (n_179), .Q (n_2205));
  AN21X1 g50114(.A (n_1423), .B (n_1422), .C (n_1), .Q (n_2204));
  AN21X1 g50111(.A (n_1421), .B (n_1420), .C (n_179), .Q (n_2203));
  AN21X1 g50110(.A (n_1419), .B (n_1418), .C (n_1), .Q (n_2202));
  AN21X1 g50104(.A (n_8321), .B (n_1416), .C (n_1), .Q (n_2201));
  AN21X1 g50094(.A (n_1415), .B (n_1414), .C (n_1), .Q (n_2200));
  AN21X1 g50082(.A (n_1413), .B (n_1412), .C (n_1), .Q (n_2199));
  AN21X1 g50105(.A (n_1411), .B (n_1410), .C (n_1), .Q (n_2198));
  AN21X1 g50097(.A (n_1409), .B (n_1408), .C (n_1), .Q (n_2197));
  AN21X1 g50083(.A (n_1407), .B (n_1406), .C (n_180), .Q (n_2196));
  AN21X1 g50072(.A (n_1405), .B (n_1404), .C (n_1), .Q (n_2195));
  NO2X1 g50192(.A (n_1403), .B (n_179), .Q (n_2194));
  AN21X1 g50106(.A (n_1402), .B (n_1401), .C (n_1), .Q (n_2193));
  AN21X1 g50095(.A (n_1400), .B (n_1399), .C (n_1), .Q (n_2192));
  AN21X1 g50084(.A (n_1398), .B (n_1397), .C (n_1), .Q (n_2191));
  AN21X1 g50074(.A (n_1396), .B (n_1395), .C (n_1), .Q (n_2190));
  AN21X1 g50096(.A (n_1394), .B (n_1393), .C (n_1), .Q (n_2189));
  AN21X1 g50085(.A (n_1392), .B (n_1391), .C (n_1), .Q (n_2188));
  AN21X1 g50075(.A (n_1390), .B (n_1389), .C (n_1), .Q (n_2187));
  AN21X1 g50062(.A (n_1388), .B (n_1387), .C (n_180), .Q (n_2186));
  AN21X1 g50098(.A (n_1386), .B (n_1385), .C (n_1), .Q (n_2185));
  AN21X1 g50086(.A (n_1384), .B (n_1383), .C (n_180), .Q (n_2184));
  NO2X1 g50190(.A (n_1382), .B (n_179), .Q (n_2183));
  AN21X1 g50076(.A (n_1381), .B (n_1380), .C (n_1), .Q (n_2182));
  AN21X1 g50063(.A (n_1379), .B (n_1378), .C (n_180), .Q (n_2181));
  AN21X1 g50087(.A (n_1377), .B (n_1376), .C (n_180), .Q (n_2180));
  AN21X1 g50073(.A (n_1375), .B (n_1374), .C (n_1), .Q (n_2179));
  AN21X1 g50064(.A (n_1373), .B (n_1372), .C (n_180), .Q (n_2178));
  AN21X1 g50057(.A (n_8323), .B (n_1370), .C (n_180), .Q (n_2177));
  AN21X1 g50067(.A (n_1369), .B (n_1368), .C (n_1), .Q (n_2176));
  AN21X1 g50059(.A (n_1367), .B (n_1366), .C (n_180), .Q (n_2175));
  AN21X1 g50056(.A (n_1365), .B (n_1364), .C (n_180), .Q (n_2174));
  AN21X1 g50050(.A (n_1363), .B (n_1362), .C (n_180), .Q (n_2173));
  NO2X1 g50186(.A (n_1361), .B (n_180), .Q (n_2172));
  AN21X1 g50060(.A (n_1360), .B (n_1359), .C (n_180), .Q (n_2171));
  NO2X1 g50053(.A (n_1358), .B (n_179), .Q (n_2170));
  AN21X1 g50048(.A (n_1357), .B (n_1356), .C (n_180), .Q (n_2169));
  AN21X1 g50049(.A (n_8661), .B (n_1354), .C (n_180), .Q (n_2168));
  NO2X1 g50170(.A (n_1353), .B (n_179), .Q (n_2167));
  NO2X1 g50161(.A (n_1352), .B (n_180), .Q (n_2166));
  NO2X1 g50162(.A (n_1351), .B (n_179), .Q (n_2165));
  NO2X1 g50157(.A (n_1350), .B (n_179), .Q (n_2164));
  AN21X1 g91868(.A (n_1349), .B (n_1348), .C (n_1), .Q (n_2163));
  AN21X1 g91869(.A (n_1347), .B (n_1346), .C (n_1), .Q (n_2162));
  AN21X1 g91870(.A (n_1345), .B (n_1344), .C (n_1), .Q (n_2161));
  AN21X1 g91871(.A (n_1343), .B (n_1342), .C (n_1), .Q (n_2160));
  AN21X1 g91872(.A (n_1341), .B (n_1340), .C (n_180), .Q (n_2159));
  AN21X1 g91873(.A (n_1339), .B (n_1338), .C (n_180), .Q (n_2158));
  AN21X1 g91874(.A (n_1337), .B (n_1336), .C (n_179), .Q (n_2157));
  AN21X1 g91875(.A (n_1335), .B (n_1334), .C (n_179), .Q (n_2156));
  AN21X1 g91876(.A (n_1333), .B (n_1332), .C (n_1), .Q (n_2155));
  AN21X1 g91877(.A (n_1331), .B (n_1330), .C (n_180), .Q (n_2154));
  AN21X1 g91878(.A (n_1329), .B (n_1328), .C (n_1), .Q (n_2153));
  AN21X1 g91879(.A (n_1327), .B (n_1326), .C (n_1), .Q (n_2152));
  AN21X1 g91880(.A (n_1325), .B (n_1324), .C (n_179), .Q (n_2151));
  AN21X1 g91881(.A (n_1323), .B (n_1322), .C (n_1), .Q (n_2150));
  AN21X1 g91882(.A (n_1321), .B (n_1320), .C (n_180), .Q (n_2149));
  AN21X1 g91883(.A (n_1319), .B (n_1318), .C (n_180), .Q (n_2148));
  AN21X1 g91884(.A (n_1317), .B (n_1316), .C (n_180), .Q (n_2147));
  AN21X1 g91885(.A (n_1315), .B (n_1314), .C (n_1), .Q (n_2146));
  AN21X1 g91886(.A (n_1313), .B (n_1312), .C (n_1), .Q (n_2145));
  AN21X1 g91887(.A (n_1311), .B (n_1310), .C (n_180), .Q (n_2144));
  AN21X1 g91888(.A (n_1309), .B (n_1308), .C (n_180), .Q (n_2143));
  AN21X1 g91889(.A (n_1307), .B (n_1306), .C (n_1), .Q (n_2142));
  AN21X1 g91890(.A (n_1305), .B (n_1304), .C (n_1), .Q (n_2141));
  AN21X1 g91891(.A (n_1303), .B (n_1302), .C (n_1), .Q (n_2140));
  AN21X1 g91892(.A (n_1301), .B (n_1300), .C (n_1), .Q (n_2139));
  AN21X1 g91893(.A (n_1299), .B (n_1298), .C (n_1), .Q (n_2138));
  AN21X1 g91894(.A (n_1297), .B (n_1296), .C (n_1), .Q (n_2137));
  AN21X1 g91895(.A (n_1295), .B (n_1294), .C (n_1), .Q (n_2136));
  AN21X1 g91896(.A (n_1293), .B (n_1292), .C (n_1), .Q (n_2135));
  AN21X1 g91897(.A (n_1291), .B (n_1290), .C (n_1), .Q (n_2134));
  AND2X1 g91898(.A (n_7380), .B (n_181), .Q (n_2133));
  AND2X1 g91899(.A (n_7388), .B (n_181), .Q (n_2132));
  AND2X1 g91900(.A (n_7385), .B (n_181), .Q (n_2131));
  AND2X1 g91901(.A (n_7384), .B (n_181), .Q (n_2130));
  AND2X1 g91902(.A (n_8571), .B (n_181), .Q (n_2129));
  NO2X1 g91903(.A (n_1447), .B (n_1), .Q (n_2128));
  NO2X1 g50198(.A (n_1289), .B (n_1), .Q (n_2127));
  NO2X1 g50151(.A (n_1288), .B (n_179), .Q (n_2126));
  NO2X1 g50165(.A (n_1287), .B (n_180), .Q (n_2125));
  NO2X1 g50155(.A (n_1286), .B (n_180), .Q (n_2124));
  NO2X1 g50152(.A (n_1285), .B (n_1), .Q (n_2123));
  NO2X1 g50148(.A (n_1284), .B (n_180), .Q (n_2122));
  NO2X1 g50142(.A (n_1283), .B (n_1), .Q (n_2121));
  NO2X1 g50143(.A (n_1282), .B (n_179), .Q (n_2120));
  NO2X1 g50137(.A (n_1281), .B (n_179), .Q (n_2119));
  NO2X1 g50129(.A (n_1280), .B (n_179), .Q (n_2118));
  NO2X1 g50124(.A (n_1279), .B (n_179), .Q (n_2117));
  NO2X1 g50196(.A (n_1278), .B (n_179), .Q (n_2116));
  NO2X1 g50139(.A (n_1277), .B (n_179), .Q (n_2115));
  NO2X1 g50130(.A (n_1276), .B (n_1), .Q (n_2114));
  NO2X1 g50138(.A (n_1275), .B (n_180), .Q (n_2113));
  NO2X1 g50131(.A (n_1274), .B (n_1), .Q (n_2112));
  NO2X1 g50136(.A (n_1273), .B (n_179), .Q (n_2111));
  NO2X1 g50132(.A (n_1272), .B (n_1), .Q (n_2110));
  NO2X1 g50125(.A (n_1271), .B (n_179), .Q (n_2109));
  NO2X1 g50121(.A (n_1270), .B (n_1), .Q (n_2108));
  NO2X1 g50120(.A (n_1269), .B (n_1), .Q (n_2107));
  NO2X1 g50117(.A (n_1268), .B (n_179), .Q (n_2106));
  NO2X1 g50193(.A (n_1267), .B (n_179), .Q (n_2105));
  NO2X1 g50115(.A (n_1266), .B (n_1), .Q (n_2104));
  AN21X1 g50113(.A (n_8327), .B (n_1264), .C (n_1), .Q (n_2103));
  NO2X1 g50112(.A (n_1263), .B (n_179), .Q (n_2102));
  AN21X1 g50107(.A (n_8329), .B (n_1261), .C (n_180), .Q (n_2101));
  NO2X1 g50100(.A (n_1260), .B (n_1), .Q (n_2100));
  AN21X1 g50093(.A (n_8331), .B (n_1258), .C (n_1), .Q (n_2099));
  AN21X1 g50108(.A (n_1257), .B (n_1256), .C (n_180), .Q (n_2098));
  NO2X1 g50103(.A (n_8576), .B (n_179), .Q (n_2097));
  AN21X1 g50090(.A (n_1254), .B (n_1253), .C (n_180), .Q (n_2096));
  NO2X1 g50079(.A (n_8577), .B (n_1), .Q (n_2095));
  NO2X1 g50188(.A (n_1251), .B (n_179), .Q (n_2094));
  AN21X1 g50109(.A (n_1250), .B (n_1249), .C (n_1), .Q (n_2093));
  NO2X1 g50101(.A (n_8578), .B (n_1), .Q (n_2092));
  AN21X1 g50088(.A (n_1247), .B (n_1246), .C (n_180), .Q (n_2091));
  NO2X1 g50081(.A (n_8579), .B (n_1), .Q (n_2090));
  NO2X1 g50102(.A (n_8687), .B (n_179), .Q (n_2089));
  AN21X1 g50089(.A (n_1243), .B (n_1242), .C (n_180), .Q (n_2088));
  NO2X1 g50080(.A (n_8688), .B (n_179), .Q (n_2087));
  AN21X1 g50068(.A (n_1240), .B (n_1239), .C (n_180), .Q (n_2086));
  NO2X1 g50099(.A (n_8689), .B (n_179), .Q (n_2085));
  AN21X1 g50091(.A (n_1237), .B (n_1236), .C (n_180), .Q (n_2084));
  NO2X1 g50187(.A (n_1235), .B (n_1), .Q (n_2083));
  NO2X1 g50077(.A (n_8690), .B (n_179), .Q (n_2082));
  AN21X1 g50070(.A (n_1233), .B (n_1232), .C (n_1), .Q (n_2081));
  AN21X1 g50092(.A (n_1231), .B (n_1230), .C (n_180), .Q (n_2080));
  NO2X1 g50078(.A (n_1229), .B (n_179), .Q (n_2079));
  AN21X1 g50069(.A (n_8333), .B (n_1227), .C (n_180), .Q (n_2078));
  NO2X1 g50061(.A (n_8691), .B (n_179), .Q (n_2077));
  NO2X1 g50071(.A (n_8692), .B (n_179), .Q (n_2076));
  AN21X1 g50066(.A (n_1224), .B (n_1223), .C (n_1), .Q (n_2075));
  NO2X1 g50058(.A (n_1222), .B (n_179), .Q (n_2074));
  AN21X1 g50054(.A (n_1221), .B (n_1220), .C (n_1), .Q (n_2073));
  NO2X1 g50184(.A (n_1219), .B (n_180), .Q (n_2072));
  AN21X1 g50065(.A (n_8335), .B (n_1217), .C (n_180), .Q (n_2071));
  NO2X1 g50055(.A (n_1216), .B (n_179), .Q (n_2070));
  AN21X1 g50052(.A (n_8337), .B (n_1214), .C (n_1), .Q (n_2069));
  AN21X1 g50051(.A (n_8339), .B (n_1212), .C (n_180), .Q (n_2068));
  NO2X1 g50164(.A (n_1211), .B (n_179), .Q (n_2067));
  NO2X1 g50159(.A (n_1210), .B (n_1), .Q (n_2066));
  NO2X1 g50160(.A (n_1209), .B (n_179), .Q (n_2065));
  NO2X1 g50156(.A (n_1208), .B (n_179), .Q (n_2064));
  NO2X1 g91904(.A (n_1207), .B (n_179), .Q (n_2063));
  NO2X1 g91905(.A (n_1206), .B (n_179), .Q (n_2062));
  AND2X1 g91906(.A (n_6233), .B (n_181), .Q (n_2061));
  AND2X1 g91907(.A (n_7635), .B (n_181), .Q (n_2060));
  AND2X1 g91908(.A (n_6234), .B (n_181), .Q (n_2059));
  AND2X1 g91909(.A (n_7632), .B (n_181), .Q (n_2058));
  NO2X1 g50354(.A (n_1205), .B (n_179), .Q (n_2057));
  AO211X1 g50351(.A (n_8340), .B (n_6256), .C (reset_internal_39074),
       .D (n_1203), .Q (n_2056));
  NO2X1 g50263(.A (n_1202), .B (n_179), .Q (n_2055));
  NO2X1 g50414(.A (n_1201), .B (n_179), .Q (n_2054));
  NO2X1 g50411(.A (n_1200), .B (n_179), .Q (n_2053));
  NO2X1 g50415(.A (n_1199), .B (n_179), .Q (n_2052));
  NO2X1 g50417(.A (n_1198), .B (n_179), .Q (n_2051));
  NO2X1 g50416(.A (n_1197), .B (n_179), .Q (n_2050));
  NO2X1 g50418(.A (n_1196), .B (n_179), .Q (n_2049));
  NO2X1 g50422(.A (n_1195), .B (n_179), .Q (n_2048));
  NO2X1 g50419(.A (n_1194), .B (n_179), .Q (n_2047));
  NO2X1 g50431(.A (n_1193), .B (n_179), .Q (n_2046));
  NO2X1 g50420(.A (n_1192), .B (n_179), .Q (n_2045));
  NO2X1 g50264(.A (n_1191), .B (n_179), .Q (n_2044));
  NO2X1 g50424(.A (n_1190), .B (n_179), .Q (n_2043));
  NO2X1 g50421(.A (n_1189), .B (n_179), .Q (n_2042));
  NO2X1 g50412(.A (n_1188), .B (n_179), .Q (n_2041));
  NO2X1 g50413(.A (n_1187), .B (n_179), .Q (n_2040));
  NO2X1 g50423(.A (n_1186), .B (n_179), .Q (n_2039));
  NO2X1 g50425(.A (n_1185), .B (n_179), .Q (n_2038));
  NO2X1 g50426(.A (n_1184), .B (n_179), .Q (n_2037));
  NO2X1 g50410(.A (n_1183), .B (n_179), .Q (n_2036));
  NO2X1 g50409(.A (n_1182), .B (n_179), .Q (n_2035));
  NO2X1 g50427(.A (n_1181), .B (n_179), .Q (n_2034));
  NO2X1 g50408(.A (n_1180), .B (n_179), .Q (n_2033));
  NO2X1 g50428(.A (n_1179), .B (n_179), .Q (n_2032));
  NO2X1 g50429(.A (n_1178), .B (n_179), .Q (n_2031));
  NO2X1 g50407(.A (n_1177), .B (n_179), .Q (n_2030));
  NO2X1 g50430(.A (n_1176), .B (n_179), .Q (n_2029));
  NO2X1 g50406(.A (n_1175), .B (n_179), .Q (n_2028));
  NO2X1 g50405(.A (n_1174), .B (n_179), .Q (n_2027));
  NO2X1 g50432(.A (n_1173), .B (n_179), .Q (n_2026));
  NO2X1 g50434(.A (n_1172), .B (n_179), .Q (n_2025));
  NO2X1 g50433(.A (n_1171), .B (n_179), .Q (n_2024));
  NO2X1 g91910(.A (n_1207), .B (n_1), .Q (n_2023));
  AND2X1 g91911(.A (n_7394), .B (n_181), .Q (n_2022));
  AND2X1 g91912(.A (n_7391), .B (n_181), .Q (n_2021));
  AND2X1 g91913(.A (n_7378), .B (n_181), .Q (n_2020));
  AND2X1 g91914(.A (n_6233), .B (n_181), .Q (n_2019));
  AND2X1 g91915(.A (n_7632), .B (n_181), .Q (n_2018));
  AND2X1 g91916(.A (n_6232), .B (n_181), .Q (n_2017));
  AND2X1 g91917(.A (n_6237), .B (n_181), .Q (n_2016));
  NO2X1 g91918(.A (n_1447), .B (n_1), .Q (n_2015));
  AND2X1 g91919(.A (n_7397), .B (n_181), .Q (n_2014));
  NO2X1 g91920(.A (n_1170), .B (n_179), .Q (n_2013));
  NO3X1 g91921(.A (n_1169), .B (flush_37557), .C (n_180), .Q (n_2012));
  NO3X1 g91922(.A (take_trap_39229), .B (n_1018), .C (n_180), .Q
       (n_2011));
  NO2X1 g47906(.A (n_1167), .B (n_1), .Q (n_2010));
  NO2X1 g48409(.A (n_1164), .B (n_179), .Q (n_2009));
  NO2X1 g49046(.A (n_1159), .B (n_179), .Q (n_2008));
  NO2X1 g49077(.A (n_1157), .B (n_179), .Q (n_2007));
  NO2X1 g48346(.A (n_1155), .B (n_1), .Q (n_2006));
  NO2X1 g49170(.A (n_1154), .B (n_180), .Q (n_2005));
  NO2X1 g48315(.A (n_1153), .B (n_179), .Q (n_2004));
  NO2X1 g49653(.A (n_8355), .B (n_179), .Q (n_2003));
  NO2X1 g49541(.A (n_1151), .B (n_179), .Q (n_2002));
  NO2X1 g49583(.A (n_1150), .B (n_180), .Q (n_2001));
  NO2X1 g49521(.A (n_1149), .B (n_180), .Q (n_2000));
  NO2X1 g49584(.A (n_1148), .B (n_180), .Q (n_1999));
  NO2X1 g49108(.A (n_1147), .B (n_179), .Q (n_1998));
  NO2X1 g49522(.A (n_1146), .B (n_180), .Q (n_1997));
  NO2X1 g49109(.A (n_1144), .B (n_179), .Q (n_1996));
  NO2X1 g49171(.A (n_1143), .B (n_180), .Q (n_1995));
  NO2X1 g47907(.A (n_1167), .B (n_1), .Q (n_1994));
  NO2X1 g48412(.A (n_1164), .B (n_179), .Q (n_1993));
  NO2X1 g49078(.A (n_1157), .B (n_180), .Q (n_1992));
  NO2X1 g48347(.A (n_1155), .B (n_1), .Q (n_1991));
  NO2X1 g49172(.A (n_1154), .B (n_180), .Q (n_1990));
  NO2X1 g48316(.A (n_1153), .B (n_180), .Q (n_1989));
  NO2X1 g49654(.A (n_8355), .B (n_180), .Q (n_1988));
  NO2X1 g49585(.A (n_1150), .B (n_180), .Q (n_1987));
  NO2X1 g49586(.A (n_1148), .B (n_180), .Q (n_1986));
  NO2X1 g49110(.A (n_1147), .B (n_180), .Q (n_1985));
  NO2X1 g49524(.A (n_1146), .B (n_180), .Q (n_1984));
  NO2X1 g49111(.A (n_1144), .B (n_179), .Q (n_1983));
  NO2X1 g49173(.A (n_1143), .B (n_180), .Q (n_1982));
  NO2X1 g47908(.A (n_1167), .B (n_1), .Q (n_1981));
  NO2X1 g48415(.A (n_1164), .B (n_179), .Q (n_1980));
  NO2X1 g49048(.A (n_1159), .B (n_179), .Q (n_1979));
  NO2X1 g49079(.A (n_1157), .B (n_180), .Q (n_1978));
  NO2X1 g48348(.A (n_1155), .B (n_1), .Q (n_1977));
  NO2X1 g49174(.A (n_1154), .B (n_179), .Q (n_1976));
  NO2X1 g48317(.A (n_1153), .B (n_179), .Q (n_1975));
  NO2X1 g49655(.A (n_8355), .B (n_180), .Q (n_1974));
  NO2X1 g49492(.A (n_1151), .B (n_179), .Q (n_1973));
  NO2X1 g49587(.A (n_1150), .B (n_180), .Q (n_1972));
  NO2X1 g49588(.A (n_1148), .B (n_179), .Q (n_1971));
  NO2X1 g49112(.A (n_1147), .B (n_180), .Q (n_1970));
  NO2X1 g49526(.A (n_1146), .B (n_180), .Q (n_1969));
  NO2X1 g49113(.A (n_1144), .B (n_179), .Q (n_1968));
  NO2X1 g49175(.A (n_1143), .B (n_180), .Q (n_1967));
  NO2X1 g47909(.A (n_1167), .B (n_1), .Q (n_1966));
  NO2X1 g48418(.A (n_1164), .B (n_179), .Q (n_1965));
  NO2X1 g49049(.A (n_1159), .B (n_179), .Q (n_1964));
  NO2X1 g49080(.A (n_1157), .B (n_179), .Q (n_1963));
  NO2X1 g48349(.A (n_1155), .B (n_179), .Q (n_1962));
  NO2X1 g49176(.A (n_1154), .B (n_180), .Q (n_1961));
  NO2X1 g48318(.A (n_1153), .B (n_179), .Q (n_1960));
  NO2X1 g49657(.A (n_8355), .B (n_180), .Q (n_1959));
  NO2X1 g49493(.A (n_1151), .B (n_179), .Q (n_1958));
  NO2X1 g49589(.A (n_1150), .B (n_180), .Q (n_1957));
  NO2X1 g49590(.A (n_1148), .B (n_179), .Q (n_1956));
  NO2X1 g49114(.A (n_1147), .B (n_180), .Q (n_1955));
  NO2X1 g49528(.A (n_1146), .B (n_180), .Q (n_1954));
  NO2X1 g49115(.A (n_1144), .B (n_179), .Q (n_1953));
  NO2X1 g49177(.A (n_1143), .B (n_179), .Q (n_1952));
  NO2X1 g47910(.A (n_1167), .B (n_1), .Q (n_1951));
  NO2X1 g48421(.A (n_1164), .B (n_179), .Q (n_1950));
  NO2X1 g49081(.A (n_1157), .B (n_179), .Q (n_1949));
  NO2X1 g48350(.A (n_1155), .B (n_179), .Q (n_1948));
  NO2X1 g49178(.A (n_1154), .B (n_180), .Q (n_1947));
  NO2X1 g48319(.A (n_1153), .B (n_179), .Q (n_1946));
  NO2X1 g49658(.A (n_8355), .B (n_180), .Q (n_1945));
  NO2X1 g49494(.A (n_1151), .B (n_179), .Q (n_1944));
  NO2X1 g49591(.A (n_1150), .B (n_179), .Q (n_1943));
  NO2X1 g49592(.A (n_1148), .B (n_180), .Q (n_1942));
  NO2X1 g49116(.A (n_1147), .B (n_180), .Q (n_1941));
  NO2X1 g49530(.A (n_1146), .B (n_180), .Q (n_1940));
  NO2X1 g49117(.A (n_1144), .B (n_180), .Q (n_1939));
  NO2X1 g49179(.A (n_1143), .B (n_180), .Q (n_1938));
  NO2X1 g47911(.A (n_1167), .B (n_1), .Q (n_1937));
  NO2X1 g49082(.A (n_1157), .B (n_179), .Q (n_1936));
  NO2X1 g48351(.A (n_1155), .B (n_1), .Q (n_1935));
  NO2X1 g49180(.A (n_1154), .B (n_180), .Q (n_1934));
  NO2X1 g48320(.A (n_1153), .B (n_179), .Q (n_1933));
  NO2X1 g49659(.A (n_8355), .B (n_179), .Q (n_1932));
  NO2X1 g49495(.A (n_1151), .B (n_179), .Q (n_1931));
  NO2X1 g49600(.A (n_1150), .B (n_180), .Q (n_1930));
  NO2X1 g49601(.A (n_1148), .B (n_180), .Q (n_1929));
  NO2X1 g49119(.A (n_1147), .B (n_179), .Q (n_1928));
  NO2X1 g49534(.A (n_1146), .B (n_180), .Q (n_1927));
  NO2X1 g49120(.A (n_1144), .B (n_180), .Q (n_1926));
  NO2X1 g49181(.A (n_1143), .B (n_180), .Q (n_1925));
  NO2X1 g47912(.A (n_1167), .B (n_1), .Q (n_1924));
  NO2X1 g49083(.A (n_1157), .B (n_180), .Q (n_1923));
  NO2X1 g48352(.A (n_1155), .B (n_1), .Q (n_1922));
  NO2X1 g49184(.A (n_1154), .B (n_180), .Q (n_1921));
  NO2X1 g48321(.A (n_1153), .B (n_180), .Q (n_1920));
  NO2X1 g49660(.A (n_8355), .B (n_180), .Q (n_1919));
  NO2X1 g49496(.A (n_1151), .B (n_179), .Q (n_1918));
  NO2X1 g49604(.A (n_1150), .B (n_180), .Q (n_1917));
  NO2X1 g49605(.A (n_1148), .B (n_180), .Q (n_1916));
  NO2X1 g49121(.A (n_1147), .B (n_180), .Q (n_1915));
  NO2X1 g49536(.A (n_1146), .B (n_180), .Q (n_1914));
  NO2X1 g49122(.A (n_1144), .B (n_180), .Q (n_1913));
  NO2X1 g49185(.A (n_1143), .B (n_180), .Q (n_1912));
  NO2X1 g47913(.A (n_1167), .B (n_1), .Q (n_1911));
  NO2X1 g48430(.A (n_1164), .B (n_179), .Q (n_1910));
  NO2X1 g49053(.A (n_1159), .B (n_179), .Q (n_1909));
  NO2X1 g49084(.A (n_1157), .B (n_180), .Q (n_1908));
  NO2X1 g48353(.A (n_1155), .B (n_1), .Q (n_1907));
  NO2X1 g49186(.A (n_1154), .B (n_180), .Q (n_1906));
  NO2X1 g48322(.A (n_1153), .B (n_180), .Q (n_1905));
  NO2X1 g49661(.A (n_8355), .B (n_180), .Q (n_1904));
  NO2X1 g49497(.A (n_1151), .B (n_179), .Q (n_1903));
  NO2X1 g49606(.A (n_1150), .B (n_180), .Q (n_1902));
  NO2X1 g49607(.A (n_1148), .B (n_180), .Q (n_1901));
  NO2X1 g49123(.A (n_1147), .B (n_179), .Q (n_1900));
  NO2X1 g49539(.A (n_1146), .B (n_180), .Q (n_1899));
  NO2X1 g49124(.A (n_1144), .B (n_180), .Q (n_1898));
  NO2X1 g49187(.A (n_1143), .B (n_180), .Q (n_1897));
  NO2X1 g47914(.A (n_1167), .B (n_1), .Q (n_1896));
  NO2X1 g48433(.A (n_1164), .B (n_179), .Q (n_1895));
  NO2X1 g49085(.A (n_1157), .B (n_180), .Q (n_1894));
  NO2X1 g48354(.A (n_1155), .B (n_1), .Q (n_1893));
  NO2X1 g49188(.A (n_1154), .B (n_180), .Q (n_1892));
  NO2X1 g48323(.A (n_1153), .B (n_180), .Q (n_1891));
  NO2X1 g49662(.A (n_8355), .B (n_179), .Q (n_1890));
  NO2X1 g49608(.A (n_1150), .B (n_180), .Q (n_1889));
  NO2X1 g49609(.A (n_1148), .B (n_179), .Q (n_1888));
  NO2X1 g49125(.A (n_1147), .B (n_180), .Q (n_1887));
  NO2X1 g49490(.A (n_1146), .B (n_180), .Q (n_1886));
  NO2X1 g49126(.A (n_1144), .B (n_180), .Q (n_1885));
  NO2X1 g49189(.A (n_1143), .B (n_180), .Q (n_1884));
  NO2X1 g47915(.A (n_1167), .B (n_1), .Q (n_1883));
  NO2X1 g48436(.A (n_1164), .B (n_179), .Q (n_1882));
  NO2X1 g49086(.A (n_1157), .B (n_179), .Q (n_1881));
  NO2X1 g48355(.A (n_1155), .B (n_1), .Q (n_1880));
  NO2X1 g49190(.A (n_1154), .B (n_180), .Q (n_1879));
  NO2X1 g48324(.A (n_1153), .B (n_180), .Q (n_1878));
  NO2X1 g49663(.A (n_8355), .B (n_180), .Q (n_1877));
  NO2X1 g49499(.A (n_1151), .B (n_179), .Q (n_1876));
  NO2X1 g49610(.A (n_1150), .B (n_180), .Q (n_1875));
  NO2X1 g49611(.A (n_1148), .B (n_180), .Q (n_1874));
  NO2X1 g49127(.A (n_1147), .B (n_180), .Q (n_1873));
  NO2X1 g49543(.A (n_1146), .B (n_179), .Q (n_1872));
  NO2X1 g49128(.A (n_1144), .B (n_180), .Q (n_1871));
  NO2X1 g49191(.A (n_1143), .B (n_179), .Q (n_1870));
  NO2X1 g47916(.A (n_1167), .B (n_1), .Q (n_1869));
  NO2X1 g48439(.A (n_1164), .B (n_179), .Q (n_1868));
  NO2X1 g49087(.A (n_1157), .B (n_180), .Q (n_1867));
  NO2X1 g48356(.A (n_1155), .B (n_1), .Q (n_1866));
  NO2X1 g49192(.A (n_1154), .B (n_180), .Q (n_1865));
  NO2X1 g48325(.A (n_1153), .B (n_180), .Q (n_1864));
  NO2X1 g49664(.A (n_8355), .B (n_179), .Q (n_1863));
  NO2X1 g49500(.A (n_1151), .B (n_179), .Q (n_1862));
  NO2X1 g49612(.A (n_1150), .B (n_180), .Q (n_1861));
  NO2X1 g49613(.A (n_1148), .B (n_179), .Q (n_1860));
  NO2X1 g49130(.A (n_1147), .B (n_180), .Q (n_1859));
  NO2X1 g49545(.A (n_1146), .B (n_179), .Q (n_1858));
  NO2X1 g49131(.A (n_1144), .B (n_180), .Q (n_1857));
  NO2X1 g49193(.A (n_1143), .B (n_179), .Q (n_1856));
  NO2X1 g47917(.A (n_1167), .B (n_1), .Q (n_1855));
  NO2X1 g49088(.A (n_1157), .B (n_180), .Q (n_1854));
  NO2X1 g48357(.A (n_1155), .B (n_1), .Q (n_1853));
  NO2X1 g49194(.A (n_1154), .B (n_179), .Q (n_1852));
  NO2X1 g48326(.A (n_1153), .B (n_180), .Q (n_1851));
  NO2X1 g49665(.A (n_8355), .B (n_180), .Q (n_1850));
  NO2X1 g49614(.A (n_1150), .B (n_180), .Q (n_1849));
  NO2X1 g49615(.A (n_1148), .B (n_180), .Q (n_1848));
  NO2X1 g49132(.A (n_1147), .B (n_179), .Q (n_1847));
  NO2X1 g49548(.A (n_1146), .B (n_180), .Q (n_1846));
  NO2X1 g49133(.A (n_1144), .B (n_179), .Q (n_1845));
  NO2X1 g49195(.A (n_1143), .B (n_179), .Q (n_1844));
  NO2X1 g47918(.A (n_1167), .B (n_1), .Q (n_1843));
  NO2X1 g49089(.A (n_1157), .B (n_180), .Q (n_1842));
  NO2X1 g48358(.A (n_1155), .B (n_1), .Q (n_1841));
  NO2X1 g49197(.A (n_1154), .B (n_180), .Q (n_1840));
  NO2X1 g48327(.A (n_1153), .B (n_179), .Q (n_1839));
  NO2X1 g49666(.A (n_8355), .B (n_179), .Q (n_1838));
  NO2X1 g49502(.A (n_1151), .B (n_179), .Q (n_1837));
  NO2X1 g49617(.A (n_1150), .B (n_179), .Q (n_1836));
  NO2X1 g49618(.A (n_1148), .B (n_179), .Q (n_1835));
  NO2X1 g49135(.A (n_1147), .B (n_179), .Q (n_1834));
  NO2X1 g49551(.A (n_1146), .B (n_180), .Q (n_1833));
  NO2X1 g49136(.A (n_1144), .B (n_180), .Q (n_1832));
  NO2X1 g49198(.A (n_1143), .B (n_180), .Q (n_1831));
  NO2X1 g47919(.A (n_1167), .B (n_1), .Q (n_1830));
  NO2X1 g48448(.A (n_1164), .B (n_179), .Q (n_1829));
  NO2X1 g49059(.A (n_1159), .B (n_179), .Q (n_1828));
  NO2X1 g49090(.A (n_1157), .B (n_179), .Q (n_1827));
  NO2X1 g48359(.A (n_1155), .B (n_1), .Q (n_1826));
  NO2X1 g49199(.A (n_1154), .B (n_180), .Q (n_1825));
  NO2X1 g48328(.A (n_1153), .B (n_180), .Q (n_1824));
  NO2X1 g49667(.A (n_8355), .B (n_180), .Q (n_1823));
  NO2X1 g49620(.A (n_1150), .B (n_179), .Q (n_1822));
  NO2X1 g49621(.A (n_1148), .B (n_180), .Q (n_1821));
  NO2X1 g49137(.A (n_1147), .B (n_179), .Q (n_1820));
  NO2X1 g49553(.A (n_1146), .B (n_180), .Q (n_1819));
  NO2X1 g49138(.A (n_1144), .B (n_179), .Q (n_1818));
  NO2X1 g49200(.A (n_1143), .B (n_180), .Q (n_1817));
  NO2X1 g47920(.A (n_1167), .B (n_179), .Q (n_1816));
  NO2X1 g48451(.A (n_1164), .B (n_179), .Q (n_1815));
  NO2X1 g49091(.A (n_1157), .B (n_180), .Q (n_1814));
  NO2X1 g48360(.A (n_1155), .B (n_1), .Q (n_1813));
  NO2X1 g49201(.A (n_1154), .B (n_180), .Q (n_1812));
  NO2X1 g48329(.A (n_1153), .B (n_180), .Q (n_1811));
  NO2X1 g49669(.A (n_8355), .B (n_180), .Q (n_1810));
  NO2X1 g49622(.A (n_1150), .B (n_180), .Q (n_1809));
  NO2X1 g49623(.A (n_1148), .B (n_180), .Q (n_1808));
  NO2X1 g49139(.A (n_1147), .B (n_180), .Q (n_1807));
  NO2X1 g49556(.A (n_1146), .B (n_180), .Q (n_1806));
  NO2X1 g49140(.A (n_1144), .B (n_179), .Q (n_1805));
  NO2X1 g49202(.A (n_1143), .B (n_179), .Q (n_1804));
  NO2X1 g47921(.A (n_1167), .B (n_179), .Q (n_1803));
  NO2X1 g49061(.A (n_1159), .B (n_179), .Q (n_1802));
  NO2X1 g49092(.A (n_1157), .B (n_180), .Q (n_1801));
  NO2X1 g48361(.A (n_1155), .B (n_1), .Q (n_1800));
  NO2X1 g49203(.A (n_1154), .B (n_180), .Q (n_1799));
  NO2X1 g48330(.A (n_1153), .B (n_180), .Q (n_1798));
  NO2X1 g49670(.A (n_8355), .B (n_180), .Q (n_1797));
  NO2X1 g49505(.A (n_1151), .B (n_179), .Q (n_1796));
  NO2X1 g49624(.A (n_1150), .B (n_180), .Q (n_1795));
  NO2X1 g49645(.A (n_1148), .B (n_179), .Q (n_1794));
  NO2X1 g49142(.A (n_1147), .B (n_180), .Q (n_1793));
  NO2X1 g49558(.A (n_1146), .B (n_179), .Q (n_1792));
  NO2X1 g49143(.A (n_1144), .B (n_180), .Q (n_1791));
  NO2X1 g49204(.A (n_1143), .B (n_179), .Q (n_1790));
  NO2X1 g47922(.A (n_1167), .B (n_179), .Q (n_1789));
  NO2X1 g49093(.A (n_1157), .B (n_180), .Q (n_1788));
  NO2X1 g48362(.A (n_1155), .B (n_1), .Q (n_1787));
  NO2X1 g49205(.A (n_1154), .B (n_179), .Q (n_1786));
  NO2X1 g48331(.A (n_1153), .B (n_179), .Q (n_1785));
  NO2X1 g49671(.A (n_8355), .B (n_179), .Q (n_1784));
  NO2X1 g49506(.A (n_1151), .B (n_179), .Q (n_1783));
  NO2X1 g49625(.A (n_1150), .B (n_180), .Q (n_1782));
  NO2X1 g49629(.A (n_1148), .B (n_179), .Q (n_1781));
  NO2X1 g49144(.A (n_1147), .B (n_179), .Q (n_1780));
  NO2X1 g49560(.A (n_1146), .B (n_180), .Q (n_1779));
  NO2X1 g49145(.A (n_1144), .B (n_179), .Q (n_1778));
  NO2X1 g49206(.A (n_1143), .B (n_180), .Q (n_1777));
  NO2X1 g47923(.A (n_1167), .B (n_179), .Q (n_1776));
  NO2X1 g48460(.A (n_1164), .B (n_179), .Q (n_1775));
  NO2X1 g49094(.A (n_1157), .B (n_180), .Q (n_1774));
  NO2X1 g48363(.A (n_1155), .B (n_1), .Q (n_1773));
  NO2X1 g49207(.A (n_1154), .B (n_180), .Q (n_1772));
  NO2X1 g48332(.A (n_1153), .B (n_180), .Q (n_1771));
  NO2X1 g49672(.A (n_8355), .B (n_179), .Q (n_1770));
  NO2X1 g49507(.A (n_1151), .B (n_179), .Q (n_1769));
  NO2X1 g49626(.A (n_1150), .B (n_180), .Q (n_1768));
  NO2X1 g49616(.A (n_1148), .B (n_180), .Q (n_1767));
  NO2X1 g49147(.A (n_1147), .B (n_179), .Q (n_1766));
  NO2X1 g49546(.A (n_1146), .B (n_180), .Q (n_1765));
  NO2X1 g49148(.A (n_1144), .B (n_180), .Q (n_1764));
  NO2X1 g49208(.A (n_1143), .B (n_180), .Q (n_1763));
  NO2X1 g47924(.A (n_1167), .B (n_1), .Q (n_1762));
  NO2X1 g48463(.A (n_1164), .B (n_179), .Q (n_1761));
  NO2X1 g49064(.A (n_1159), .B (n_179), .Q (n_1760));
  NO2X1 g49095(.A (n_1157), .B (n_180), .Q (n_1759));
  NO2X1 g48364(.A (n_1155), .B (n_1), .Q (n_1758));
  NO2X1 g49209(.A (n_1154), .B (n_179), .Q (n_1757));
  NO2X1 g48333(.A (n_1153), .B (n_179), .Q (n_1756));
  NO2X1 g49673(.A (n_8355), .B (n_179), .Q (n_1755));
  NO2X1 g49508(.A (n_1151), .B (n_179), .Q (n_1754));
  NO2X1 g49628(.A (n_1150), .B (n_179), .Q (n_1753));
  NO2X1 g49602(.A (n_1148), .B (n_180), .Q (n_1752));
  NO2X1 g49150(.A (n_1147), .B (n_179), .Q (n_1751));
  NO2X1 g49531(.A (n_1146), .B (n_179), .Q (n_1750));
  NO2X1 g49151(.A (n_1144), .B (n_179), .Q (n_1749));
  NO2X1 g49210(.A (n_1143), .B (n_180), .Q (n_1748));
  NO2X1 g47925(.A (n_1167), .B (n_1), .Q (n_1747));
  NO2X1 g49065(.A (n_1159), .B (n_179), .Q (n_1746));
  NO2X1 g49096(.A (n_1157), .B (n_180), .Q (n_1745));
  NO2X1 g48365(.A (n_1155), .B (n_1), .Q (n_1744));
  NO2X1 g49211(.A (n_1154), .B (n_180), .Q (n_1743));
  NO2X1 g48334(.A (n_1153), .B (n_180), .Q (n_1742));
  NO2X1 g49674(.A (n_8355), .B (n_180), .Q (n_1741));
  NO2X1 g49630(.A (n_1150), .B (n_180), .Q (n_1740));
  NO2X1 g49635(.A (n_1148), .B (n_180), .Q (n_1739));
  NO2X1 g49152(.A (n_1147), .B (n_180), .Q (n_1738));
  NO2X1 g49562(.A (n_1146), .B (n_180), .Q (n_1737));
  NO2X1 g49153(.A (n_1144), .B (n_180), .Q (n_1736));
  NO2X1 g49212(.A (n_1143), .B (n_180), .Q (n_1735));
  NO2X1 g47926(.A (n_1167), .B (n_1), .Q (n_1734));
  NO2X1 g49097(.A (n_1157), .B (n_180), .Q (n_1733));
  NO2X1 g48366(.A (n_1155), .B (n_179), .Q (n_1732));
  NO2X1 g49213(.A (n_1154), .B (n_180), .Q (n_1731));
  NO2X1 g48335(.A (n_1153), .B (n_180), .Q (n_1730));
  NO2X1 g49675(.A (n_8355), .B (n_179), .Q (n_1729));
  NO2X1 g49632(.A (n_1150), .B (n_180), .Q (n_1728));
  NO2X1 g49636(.A (n_1148), .B (n_180), .Q (n_1727));
  NO2X1 g49154(.A (n_1147), .B (n_179), .Q (n_1726));
  NO2X1 g49579(.A (n_1146), .B (n_180), .Q (n_1725));
  NO2X1 g49155(.A (n_1144), .B (n_180), .Q (n_1724));
  NO2X1 g49214(.A (n_1143), .B (n_180), .Q (n_1723));
  NO2X1 g47927(.A (n_1167), .B (n_1), .Q (n_1722));
  NO2X1 g48472(.A (n_1164), .B (n_179), .Q (n_1721));
  NO2X1 g49067(.A (n_1159), .B (n_179), .Q (n_1720));
  NO2X1 g49098(.A (n_1157), .B (n_180), .Q (n_1719));
  NO2X1 g48367(.A (n_1155), .B (n_1), .Q (n_1718));
  NO2X1 g49215(.A (n_1154), .B (n_179), .Q (n_1717));
  NO2X1 g48336(.A (n_1153), .B (n_180), .Q (n_1716));
  NO2X1 g49656(.A (n_8355), .B (n_180), .Q (n_1715));
  NO2X1 g49511(.A (n_1151), .B (n_179), .Q (n_1714));
  NO2X1 g49634(.A (n_1150), .B (n_179), .Q (n_1713));
  NO2X1 g49639(.A (n_1148), .B (n_180), .Q (n_1712));
  NO2X1 g49157(.A (n_1147), .B (n_179), .Q (n_1711));
  NO2X1 g49574(.A (n_1146), .B (n_180), .Q (n_1710));
  NO2X1 g49158(.A (n_1144), .B (n_180), .Q (n_1709));
  NO2X1 g49217(.A (n_1143), .B (n_180), .Q (n_1708));
  NO2X1 g47928(.A (n_1167), .B (n_1), .Q (n_1707));
  NO2X1 g48474(.A (n_1164), .B (n_179), .Q (n_1706));
  NO2X1 g49068(.A (n_1159), .B (n_179), .Q (n_1705));
  NO2X1 g49099(.A (n_1157), .B (n_180), .Q (n_1704));
  NO2X1 g48368(.A (n_1155), .B (n_1), .Q (n_1703));
  NO2X1 g49218(.A (n_1154), .B (n_180), .Q (n_1702));
  NO2X1 g48337(.A (n_1153), .B (n_180), .Q (n_1701));
  NO2X1 g49677(.A (n_8355), .B (n_180), .Q (n_1700));
  NO2X1 g49637(.A (n_1150), .B (n_180), .Q (n_1699));
  NO2X1 g49650(.A (n_1148), .B (n_180), .Q (n_1698));
  NO2X1 g49159(.A (n_1147), .B (n_180), .Q (n_1697));
  NO2X1 g49581(.A (n_1146), .B (n_180), .Q (n_1696));
  NO2X1 g49160(.A (n_1144), .B (n_180), .Q (n_1695));
  NO2X1 g49219(.A (n_1143), .B (n_180), .Q (n_1694));
  NO2X1 g47929(.A (n_1167), .B (n_1), .Q (n_1693));
  NO2X1 g48478(.A (n_1164), .B (n_179), .Q (n_1692));
  NO2X1 g49100(.A (n_1157), .B (n_179), .Q (n_1691));
  NO2X1 g48369(.A (n_1155), .B (n_1), .Q (n_1690));
  NO2X1 g49220(.A (n_1154), .B (n_180), .Q (n_1689));
  NO2X1 g48338(.A (n_1153), .B (n_180), .Q (n_1688));
  NO2X1 g49678(.A (n_8355), .B (n_180), .Q (n_1687));
  NO2X1 g49640(.A (n_1150), .B (n_180), .Q (n_1686));
  NO2X1 g49633(.A (n_1148), .B (n_180), .Q (n_1685));
  NO2X1 g49161(.A (n_1147), .B (n_179), .Q (n_1684));
  NO2X1 g49567(.A (n_1146), .B (n_180), .Q (n_1683));
  NO2X1 g49146(.A (n_1144), .B (n_180), .Q (n_1682));
  NO2X1 g49221(.A (n_1143), .B (n_179), .Q (n_1681));
  NO2X1 g47930(.A (n_1167), .B (n_1), .Q (n_1680));
  NO2X1 g48481(.A (n_1164), .B (n_179), .Q (n_1679));
  NO2X1 g49101(.A (n_1157), .B (n_179), .Q (n_1678));
  NO2X1 g48370(.A (n_1155), .B (n_1), .Q (n_1677));
  NO2X1 g49222(.A (n_1154), .B (n_179), .Q (n_1676));
  NO2X1 g48339(.A (n_1153), .B (n_179), .Q (n_1675));
  NO2X1 g49679(.A (n_8355), .B (n_180), .Q (n_1674));
  NO2X1 g49514(.A (n_1151), .B (n_179), .Q (n_1673));
  NO2X1 g49641(.A (n_1150), .B (n_179), .Q (n_1672));
  NO2X1 g49648(.A (n_1148), .B (n_179), .Q (n_1671));
  NO2X1 g49163(.A (n_1147), .B (n_179), .Q (n_1670));
  NO2X1 g49537(.A (n_1146), .B (n_180), .Q (n_1669));
  NO2X1 g49156(.A (n_1144), .B (n_179), .Q (n_1668));
  NO2X1 g49223(.A (n_1143), .B (n_180), .Q (n_1667));
  NO2X1 g47931(.A (n_1167), .B (n_1), .Q (n_1666));
  NO2X1 g48484(.A (n_1164), .B (n_179), .Q (n_1665));
  NO2X1 g49102(.A (n_1157), .B (n_180), .Q (n_1664));
  NO2X1 g48371(.A (n_1155), .B (n_1), .Q (n_1663));
  NO2X1 g49224(.A (n_1154), .B (n_180), .Q (n_1662));
  NO2X1 g48340(.A (n_1153), .B (n_179), .Q (n_1661));
  NO2X1 g49680(.A (n_8355), .B (n_180), .Q (n_1660));
  NO2X1 g49515(.A (n_1151), .B (n_179), .Q (n_1659));
  NO2X1 g49642(.A (n_1150), .B (n_180), .Q (n_1658));
  NO2X1 g49638(.A (n_1148), .B (n_180), .Q (n_1657));
  NO2X1 g49164(.A (n_1147), .B (n_179), .Q (n_1656));
  NO2X1 g49564(.A (n_1146), .B (n_179), .Q (n_1655));
  NO2X1 g49141(.A (n_1144), .B (n_179), .Q (n_1654));
  NO2X1 g49225(.A (n_1143), .B (n_179), .Q (n_1653));
  NO2X1 g47932(.A (n_1167), .B (n_1), .Q (n_1652));
  NO2X1 g48487(.A (n_1164), .B (n_179), .Q (n_1651));
  NO2X1 g49103(.A (n_1157), .B (n_180), .Q (n_1650));
  NO2X1 g48372(.A (n_1155), .B (n_1), .Q (n_1649));
  NO2X1 g49226(.A (n_1154), .B (n_179), .Q (n_1648));
  NO2X1 g48341(.A (n_1153), .B (n_180), .Q (n_1647));
  NO2X1 g49682(.A (n_8355), .B (n_180), .Q (n_1646));
  NO2X1 g49516(.A (n_1151), .B (n_179), .Q (n_1645));
  NO2X1 g49644(.A (n_1150), .B (n_180), .Q (n_1644));
  NO2X1 g49643(.A (n_1148), .B (n_180), .Q (n_1643));
  NO2X1 g49165(.A (n_1147), .B (n_179), .Q (n_1642));
  NO2X1 g49576(.A (n_1146), .B (n_180), .Q (n_1641));
  NO2X1 g49162(.A (n_1144), .B (n_179), .Q (n_1640));
  NO2X1 g49227(.A (n_1143), .B (n_179), .Q (n_1639));
  NO2X1 g47933(.A (n_1167), .B (n_179), .Q (n_1638));
  NO2X1 g49073(.A (n_1159), .B (n_179), .Q (n_1637));
  NO2X1 g49104(.A (n_1157), .B (n_179), .Q (n_1636));
  NO2X1 g48373(.A (n_1155), .B (n_1), .Q (n_1635));
  NO2X1 g49216(.A (n_1154), .B (n_180), .Q (n_1634));
  NO2X1 g48342(.A (n_1153), .B (n_180), .Q (n_1633));
  NO2X1 g49676(.A (n_8355), .B (n_179), .Q (n_1632));
  NO2X1 g49517(.A (n_1151), .B (n_179), .Q (n_1631));
  NO2X1 g49646(.A (n_1150), .B (n_180), .Q (n_1630));
  NO2X1 g49631(.A (n_1148), .B (n_180), .Q (n_1629));
  NO2X1 g49166(.A (n_1147), .B (n_179), .Q (n_1628));
  NO2X1 g49565(.A (n_1146), .B (n_180), .Q (n_1627));
  NO2X1 g49149(.A (n_1144), .B (n_180), .Q (n_1626));
  NO2X1 g49228(.A (n_1143), .B (n_180), .Q (n_1625));
  NO2X1 g47934(.A (n_1167), .B (n_179), .Q (n_1624));
  NO2X1 g49105(.A (n_1157), .B (n_179), .Q (n_1623));
  NO2X1 g48374(.A (n_1155), .B (n_1), .Q (n_1622));
  NO2X1 g49196(.A (n_1154), .B (n_179), .Q (n_1621));
  NO2X1 g48343(.A (n_1153), .B (n_179), .Q (n_1620));
  NO2X1 g49668(.A (n_8355), .B (n_179), .Q (n_1619));
  NO2X1 g49647(.A (n_1150), .B (n_180), .Q (n_1618));
  NO2X1 g49619(.A (n_1148), .B (n_180), .Q (n_1617));
  NO2X1 g49167(.A (n_1147), .B (n_180), .Q (n_1616));
  NO2X1 g49549(.A (n_1146), .B (n_180), .Q (n_1615));
  NO2X1 g49134(.A (n_1144), .B (n_180), .Q (n_1614));
  NO2X1 g49229(.A (n_1143), .B (n_180), .Q (n_1613));
  NO2X1 g47935(.A (n_1167), .B (n_1), .Q (n_1612));
  NO2X1 g49106(.A (n_1157), .B (n_180), .Q (n_1611));
  NO2X1 g48375(.A (n_1155), .B (n_1), .Q (n_1610));
  NO2X1 g49182(.A (n_1154), .B (n_180), .Q (n_1609));
  NO2X1 g48344(.A (n_1153), .B (n_179), .Q (n_1608));
  NO2X1 g49652(.A (n_8355), .B (n_180), .Q (n_1607));
  NO2X1 g49649(.A (n_1150), .B (n_180), .Q (n_1606));
  NO2X1 g49603(.A (n_1148), .B (n_180), .Q (n_1605));
  NO2X1 g49168(.A (n_1147), .B (n_179), .Q (n_1604));
  NO2X1 g49532(.A (n_1146), .B (n_180), .Q (n_1603));
  NO2X1 g49118(.A (n_1144), .B (n_180), .Q (n_1602));
  NO2X1 g49230(.A (n_1143), .B (n_180), .Q (n_1601));
  NO2X1 g47844(.A (n_1167), .B (n_1), .Q (n_1600));
  NO2X1 g49076(.A (n_1159), .B (n_179), .Q (n_1599));
  NO2X1 g49107(.A (n_1157), .B (n_180), .Q (n_1598));
  NO2X1 g48376(.A (n_1155), .B (n_1), .Q (n_1597));
  NO2X1 g49183(.A (n_1154), .B (n_180), .Q (n_1596));
  NO2X1 g48345(.A (n_1153), .B (n_180), .Q (n_1595));
  NO2X1 g49681(.A (n_8355), .B (n_179), .Q (n_1594));
  NO2X1 g49651(.A (n_1150), .B (n_180), .Q (n_1593));
  NO2X1 g49627(.A (n_1148), .B (n_180), .Q (n_1592));
  NO2X1 g49169(.A (n_1147), .B (n_180), .Q (n_1591));
  NO2X1 g49554(.A (n_1146), .B (n_180), .Q (n_1590));
  NO2X1 g49129(.A (n_1144), .B (n_179), .Q (n_1589));
  NO2X1 g49231(.A (n_1143), .B (n_179), .Q (n_1588));
  AND2X1 g91923(.A (\instruction_address[0] ), .B (n_181), .Q (n_1587));
  OR2X1 g91924(.A (instruction[0]), .B (n_1), .Q (n_1586));
  AND2X1 g91925(.A (\instruction[10]_40063 ), .B (n_181), .Q (n_1585));
  AND2X1 g91926(.A (\instruction[11]_40312 ), .B (n_181), .Q (n_1584));
  AND2X1 g91927(.A (n_8676), .B (n_181), .Q (n_1583));
  AND2X1 g91928(.A (n_8487), .B (n_181), .Q (n_1582));
  AND2X1 g91929(.A (\instruction[14]_40189 ), .B (n_181), .Q (n_1581));
  AND2X1 g91930(.A (instruction[15]), .B (n_181), .Q (n_1580));
  AND2X1 g91931(.A (n_4643), .B (n_181), .Q (n_1579));
  AND2X1 g91932(.A (instruction[17]), .B (n_181), .Q (n_1578));
  AND2X1 g91933(.A (instruction[18]), .B (n_181), .Q (n_1577));
  AND2X1 g91934(.A (n_4640), .B (n_181), .Q (n_1576));
  OR2X1 g91935(.A (instruction[1]), .B (n_1), .Q (n_1575));
  AND2X1 g91936(.A (instruction[20]), .B (n_181), .Q (n_1574));
  AND2X1 g91937(.A (instruction[21]), .B (n_181), .Q (n_1573));
  AND2X1 g91938(.A (instruction[22]), .B (n_181), .Q (n_1572));
  AND2X1 g91939(.A (instruction[23]), .B (n_181), .Q (n_1571));
  AND2X1 g91940(.A (instruction[24]), .B (n_181), .Q (n_1570));
  AND2X1 g91941(.A (n_8485), .B (n_181), .Q (n_1569));
  AND2X1 g91942(.A (n_8486), .B (n_181), .Q (n_1568));
  AND2X1 g91943(.A (n_8480), .B (n_181), .Q (n_1567));
  AND2X1 g91944(.A (instruction[28]), .B (n_181), .Q (n_1566));
  AND2X1 g91945(.A (n_8481), .B (n_181), .Q (n_1565));
  AND2X1 g91946(.A (instruction[2]), .B (n_181), .Q (n_1564));
  AND2X1 g91947(.A (n_8484), .B (n_181), .Q (n_1563));
  AND2X1 g91948(.A (n_8482), .B (n_181), .Q (n_1562));
  AND2X1 g91949(.A (instruction[3]), .B (n_181), .Q (n_1561));
  OR2X1 g91950(.A (instruction[4]), .B (n_1), .Q (n_1560));
  AND2X1 g91951(.A (\instruction[5]_40251 ), .B (n_181), .Q (n_1559));
  AND2X1 g91952(.A (instruction[6]), .B (n_181), .Q (n_1558));
  AND2X1 g91953(.A (\instruction[7]_39642 ), .B (n_181), .Q (n_1557));
  AND2X1 g91954(.A (\instruction[8]_40127 ), .B (n_181), .Q (n_1556));
  AND2X1 g91955(.A (\instruction[9]_40095 ), .B (n_181), .Q (n_1555));
  NO2X1 g91956(.A (load_request_BAR), .B (n_179), .Q (n_1554));
  AND2X1 g91957(.A (read_request), .B (n_181), .Q (n_1553));
  NO2X1 g91958(.A (n_1135), .B (n_179), .Q (n_1552));
  NO2X1 g91959(.A (n_1134), .B (n_1), .Q (n_1551));
  NO2X1 g91960(.A (n_1133), .B (n_179), .Q (n_1550));
  NO2X1 g91961(.A (n_1132), .B (n_179), .Q (n_1549));
  NO2X1 g91962(.A (n_1131), .B (n_179), .Q (n_1548));
  NO2X1 g51538(.A (n_1130), .B (n_179), .Q (n_1547));
  NO2X1 g91963(.A (n_1129), .B (n_1), .Q (n_1546));
  NO2X1 g91964(.A (n_1128), .B (n_1), .Q (n_1545));
  NO2X1 g91965(.A (n_1127), .B (n_179), .Q (n_1544));
  NO2X1 g91966(.A (n_1126), .B (n_179), .Q (n_1543));
  NO2X1 g91967(.A (n_1125), .B (n_1), .Q (n_1542));
  NO2X1 g91968(.A (n_1124), .B (n_1), .Q (n_1541));
  NO2X1 g91969(.A (n_1123), .B (n_1), .Q (n_1540));
  NO2X1 g91970(.A (n_1122), .B (n_1), .Q (n_1539));
  NO2X1 g91971(.A (n_1121), .B (n_179), .Q (n_1538));
  NO2X1 g91972(.A (n_1120), .B (n_179), .Q (n_1537));
  NO2X1 g91973(.A (n_1119), .B (n_1), .Q (n_1536));
  NO2X1 g91974(.A (n_1118), .B (n_1), .Q (n_1535));
  NO2X1 g91975(.A (n_1117), .B (n_179), .Q (n_1534));
  NO2X1 g91976(.A (n_1116), .B (n_179), .Q (n_1533));
  NO2X1 g91977(.A (n_1115), .B (n_1), .Q (n_1532));
  NO2X1 g91978(.A (n_1114), .B (n_179), .Q (n_1531));
  NO2X1 g91979(.A (n_1113), .B (n_1), .Q (n_1530));
  NO2X1 g91980(.A (n_1112), .B (n_1), .Q (n_1529));
  NO2X1 g91981(.A (n_1111), .B (n_1), .Q (n_1528));
  NO2X1 g91982(.A (n_1110), .B (n_1), .Q (n_1527));
  NO2X1 g91983(.A (n_1109), .B (n_179), .Q (n_1526));
  NO2X1 g91984(.A (n_1108), .B (n_1), .Q (n_1525));
  NO2X1 g91985(.A (n_1107), .B (n_1), .Q (n_1524));
  NO2X1 g91986(.A (n_1106), .B (n_1), .Q (n_1523));
  AND2X1 g91987(.A (write_data[0]), .B (n_181), .Q (n_1522));
  AND2X1 g91988(.A (write_data[10]), .B (n_181), .Q (n_1521));
  AND2X1 g91989(.A (write_data[11]), .B (n_181), .Q (n_1520));
  AND2X1 g91990(.A (write_data[12]), .B (n_181), .Q (n_1519));
  AND2X1 g91991(.A (write_data[13]), .B (n_181), .Q (n_1518));
  AND2X1 g91992(.A (write_data[14]), .B (n_181), .Q (n_1517));
  AND2X1 g91993(.A (write_data[15]), .B (n_181), .Q (n_1516));
  AND2X1 g91994(.A (write_data[16]), .B (n_181), .Q (n_1515));
  AND2X1 g91995(.A (write_data[17]), .B (n_181), .Q (n_1514));
  AND2X1 g91996(.A (write_data[18]), .B (n_181), .Q (n_1513));
  AND2X1 g91997(.A (write_data[19]), .B (n_181), .Q (n_1512));
  AND2X1 g91998(.A (write_data[1]), .B (n_181), .Q (n_1511));
  AND2X1 g91999(.A (write_data[20]), .B (n_181), .Q (n_1510));
  AND2X1 g92000(.A (write_data[21]), .B (n_181), .Q (n_1509));
  AND2X1 g92001(.A (write_data[22]), .B (n_181), .Q (n_1508));
  AND2X1 g92002(.A (write_data[23]), .B (n_181), .Q (n_1507));
  AND2X1 g92003(.A (write_data[24]), .B (n_181), .Q (n_1506));
  AND2X1 g92004(.A (write_data[25]), .B (n_181), .Q (n_1505));
  AND2X1 g92005(.A (write_data[26]), .B (n_181), .Q (n_1504));
  AND2X1 g92006(.A (write_data[27]), .B (n_181), .Q (n_1503));
  AND2X1 g92007(.A (write_data[28]), .B (n_181), .Q (n_1502));
  AND2X1 g92008(.A (write_data[29]), .B (n_181), .Q (n_1501));
  AND2X1 g92009(.A (write_data[2]), .B (n_181), .Q (n_1500));
  AND2X1 g92010(.A (write_data[30]), .B (n_181), .Q (n_1499));
  AND2X1 g92011(.A (write_data[31]), .B (n_181), .Q (n_1498));
  AND2X1 g92012(.A (write_data[3]), .B (n_181), .Q (n_1497));
  AND2X1 g92013(.A (write_data[4]), .B (n_181), .Q (n_1496));
  AND2X1 g92014(.A (write_data[5]), .B (n_181), .Q (n_1495));
  AND2X1 g92015(.A (write_data[6]), .B (n_181), .Q (n_1494));
  AND2X1 g92016(.A (write_data[7]), .B (n_181), .Q (n_1493));
  AND2X1 g92017(.A (write_data[8]), .B (n_181), .Q (n_1492));
  AND2X1 g92018(.A (write_data[9]), .B (n_181), .Q (n_1491));
  AND2X1 g92019(.A (write_request), .B (n_181), .Q (n_1490));
  AND2X1 g92020(.A (n_7629), .B (n_181), .Q (n_1489));
  AND2X1 g92021(.A (n_7631), .B (n_181), .Q (n_1488));
  AND2X1 g92022(.A (n_7628), .B (n_181), .Q (n_1487));
  AND2X1 g92023(.A (n_8231), .B (n_181), .Q (n_1486));
  AND2X1 g92024(.A (n_8242), .B (n_181), .Q (n_1485));
  AND2X1 g92025(.A (n_8243), .B (n_181), .Q (n_1484));
  AND2X1 g92026(.A (n_8244), .B (n_181), .Q (n_1483));
  AND2X1 g92027(.A (n_8246), .B (n_181), .Q (n_1482));
  AND2X1 g92028(.A (n_8247), .B (n_181), .Q (n_1481));
  AND2X1 g92029(.A (n_8248), .B (n_181), .Q (n_1480));
  AND2X1 g92030(.A (n_8249), .B (n_181), .Q (n_1479));
  AND2X1 g92031(.A (n_8250), .B (n_181), .Q (n_1478));
  AND2X1 g92032(.A (n_8251), .B (n_181), .Q (n_1477));
  AND2X1 g92033(.A (n_8252), .B (n_181), .Q (n_1476));
  AND2X1 g92034(.A (n_8232), .B (n_181), .Q (n_1475));
  AND2X1 g92035(.A (n_8253), .B (n_181), .Q (n_1474));
  AND2X1 g92036(.A (n_8254), .B (n_181), .Q (n_1473));
  AND2X1 g92037(.A (n_8255), .B (n_181), .Q (n_1472));
  AND2X1 g92038(.A (n_8225), .B (n_181), .Q (n_1471));
  AND2X1 g92039(.A (n_8226), .B (n_181), .Q (n_1470));
  AND2X1 g92040(.A (n_8227), .B (n_181), .Q (n_1469));
  AND2X1 g92041(.A (n_8228), .B (n_181), .Q (n_1468));
  AND2X1 g92042(.A (n_8229), .B (n_181), .Q (n_1467));
  AND2X1 g92043(.A (n_8230), .B (n_181), .Q (n_1466));
  AND2X1 g92044(.A (n_8234), .B (n_181), .Q (n_1465));
  AND2X1 g92045(.A (n_8233), .B (n_181), .Q (n_1464));
  AND2X1 g92046(.A (n_8245), .B (n_181), .Q (n_1463));
  AND2X1 g92047(.A (n_8256), .B (n_181), .Q (n_1462));
  AND2X1 g92048(.A (n_8235), .B (n_181), .Q (n_1461));
  AND2X1 g92049(.A (n_8236), .B (n_181), .Q (n_1460));
  AND2X1 g92050(.A (n_8237), .B (n_181), .Q (n_1459));
  AND2X1 g92051(.A (n_8238), .B (n_181), .Q (n_1458));
  AND2X1 g92052(.A (n_8239), .B (n_181), .Q (n_1457));
  AND2X1 g92053(.A (n_8240), .B (n_181), .Q (n_1456));
  AND2X1 g92054(.A (n_8241), .B (n_181), .Q (n_1455));
  NO3X1 g50958(.A (n_8211), .B (n_8209), .C (n_8210), .Q (n_1454));
  MU2IX1 g92055(.S (n_8078), .IN0 (csr_mcause_code[0]), .IN1 (n_6236),
       .Q (n_1453));
  MU2IX1 g92056(.S (n_8078), .IN0 (csr_mcause_code[1]), .IN1 (n_6235),
       .Q (n_1452));
  MU2IX1 g92057(.S (n_8078), .IN0 (csr_mcause_code[2]), .IN1 (n_6233),
       .Q (n_1451));
  MU2IX1 g92058(.S (n_8078), .IN0 (csr_mcause_interrupt_flag), .IN1
       (n_7635), .Q (n_1450));
  MU2IX1 g92059(.S (n_8078), .IN0 (csr_mcause_code[3]), .IN1 (n_6234),
       .Q (n_1449));
  MU2IX1 g92060(.S (n_8078), .IN0 (csr_mcause_code[4]), .IN1 (n_7632),
       .Q (n_1448));
  INX1 g92061(.A (n_6238), .Q (n_1447));
  ON22X1 g50363(.A (n_1105), .B (csr_mcycle[0]), .C (n_6236), .D
       (n_178), .Q (n_1446));
  AN222X1 g50302(.A (n_8137), .B (n_8361), .C (n_8138), .D (n_8588), .E
       (n_7997), .F (n_8587), .Q (n_1445));
  AN222X1 g50298(.A (n_8135), .B (n_8361), .C (n_8136), .D (n_8588), .E
       (n_7996), .F (n_8587), .Q (n_1444));
  AN222X1 g50307(.A (n_8133), .B (n_8361), .C (n_8134), .D (n_8588), .E
       (n_7995), .F (n_8587), .Q (n_1443));
  AN222X1 g50303(.A (n_8131), .B (n_8361), .C (n_8132), .D (n_8588), .E
       (n_7994), .F (n_8587), .Q (n_1442));
  AN222X1 g50299(.A (n_8129), .B (n_8361), .C (n_8130), .D (n_8588), .E
       (n_7993), .F (n_8587), .Q (n_1441));
  AN222X1 g50294(.A (n_8127), .B (n_8361), .C (n_8128), .D (n_8588), .E
       (n_7992), .F (n_8587), .Q (n_1440));
  AN222X1 g50295(.A (n_8125), .B (n_8361), .C (n_8126), .D (n_8588), .E
       (n_7991), .F (n_8587), .Q (n_1439));
  AN222X1 g50290(.A (n_8361), .B (n_8123), .C (n_8124), .D (n_8588), .E
       (n_175), .F (n_7990), .Q (n_1438));
  AN222X1 g50283(.A (n_8361), .B (n_8121), .C (n_8588), .D (n_8122), .E
       (n_175), .F (n_7989), .Q (n_1437));
  AN222X1 g50276(.A (n_8361), .B (n_8119), .C (n_8588), .D (n_8120), .E
       (n_175), .F (n_7988), .Q (n_1436));
  AN222X1 g50352(.A (n_8155), .B (n_8361), .C (n_8156), .D (n_8588), .E
       (n_8006), .F (n_8587), .Q (n_1435));
  AN222X1 g50291(.A (n_8361), .B (n_8117), .C (n_8118), .D (n_8588), .E
       (n_175), .F (n_7987), .Q (n_1434));
  AN222X1 g50284(.A (n_8361), .B (n_8115), .C (n_8588), .D (n_8116), .E
       (n_175), .F (n_7986), .Q (n_1433));
  AN222X1 g50277(.A (n_8361), .B (n_8113), .C (n_8588), .D (n_8114), .E
       (n_175), .F (n_7985), .Q (n_1432));
  AN222X1 g50272(.A (n_8111), .B (n_8361), .C (n_8588), .D (n_8112), .E
       (n_175), .F (n_7984), .Q (n_1431));
  AN222X1 g50285(.A (n_8361), .B (n_8109), .C (n_8588), .D (n_8110), .E
       (n_175), .F (n_7983), .Q (n_1430));
  AN222X1 g50278(.A (n_8361), .B (n_8107), .C (n_8588), .D (n_8108), .E
       (n_175), .F (n_7982), .Q (n_1429));
  AN222X1 g50273(.A (n_8105), .B (n_8361), .C (n_8588), .D (n_8106), .E
       (n_175), .F (n_7981), .Q (n_1428));
  AN222X1 g50268(.A (n_8103), .B (n_8361), .C (n_8588), .D (n_8104), .E
       (n_175), .F (n_7980), .Q (n_1427));
  AN222X1 g50269(.A (n_8361), .B (n_8101), .C (n_8588), .D (n_8102), .E
       (n_175), .F (n_7979), .Q (n_1426));
  AN222X1 g50266(.A (n_8099), .B (n_8361), .C (n_8588), .D (n_8100), .E
       (n_175), .F (n_7978), .Q (n_1425));
  AN222X1 g50349(.A (n_8153), .B (n_8361), .C (n_8154), .D (n_8588), .E
       (n_8005), .F (n_8587), .Q (n_1424));
  NA2X1 g92062(.A (n_7977), .B (n_175), .Q (n_1423));
  AN22X1 g50560(.A (n_8097), .B (n_8361), .C (n_8098), .D (n_8588), .Q
       (n_1422));
  NA2X1 g92063(.A (n_7976), .B (n_175), .Q (n_1421));
  AN22X1 g50545(.A (n_8095), .B (n_8361), .C (n_8096), .D (n_8588), .Q
       (n_1420));
  NA2X1 g92064(.A (n_7975), .B (n_175), .Q (n_1419));
  AN22X1 g50543(.A (n_8093), .B (n_8361), .C (n_8094), .D (n_8588), .Q
       (n_1418));
  AN22X1 g50532(.A (n_8091), .B (n_8361), .C (n_8092), .D (n_8588), .Q
       (n_1416));
  NA2X1 g92066(.A (n_7973), .B (n_175), .Q (n_1415));
  AN22X1 g50516(.A (n_8089), .B (n_8361), .C (n_8090), .D (n_8588), .Q
       (n_1414));
  NA2X1 g92067(.A (n_7972), .B (n_175), .Q (n_1413));
  AN22X1 g50512(.A (n_8087), .B (n_8361), .C (n_8088), .D (n_8588), .Q
       (n_1412));
  NA2X1 g92068(.A (n_7971), .B (n_175), .Q (n_1411));
  AN22X1 g50515(.A (n_8085), .B (n_8361), .C (n_8086), .D (n_8588), .Q
       (n_1410));
  NA2X1 g92069(.A (n_7970), .B (n_175), .Q (n_1409));
  AN22X1 g50509(.A (n_8083), .B (n_8361), .C (n_8084), .D (n_8588), .Q
       (n_1408));
  NA2X1 g92070(.A (n_7969), .B (n_175), .Q (n_1407));
  AN22X1 g50488(.A (n_8081), .B (n_8361), .C (n_8082), .D (n_8588), .Q
       (n_1406));
  NA2X1 g92071(.A (n_7968), .B (n_175), .Q (n_1405));
  AN22X1 g50479(.A (n_8079), .B (n_8361), .C (n_8080), .D (n_8588), .Q
       (n_1404));
  AN222X1 g50346(.A (n_8151), .B (n_8361), .C (n_8152), .D (n_8588), .E
       (n_8004), .F (n_8587), .Q (n_1403));
  NA2X1 g92072(.A (n_7967), .B (n_175), .Q (n_1402));
  AN22X1 g50507(.A (n_8076), .B (n_8361), .C (n_8077), .D (n_8588), .Q
       (n_1401));
  NA2X1 g92073(.A (n_7966), .B (n_175), .Q (n_1400));
  AN22X1 g50485(.A (n_8074), .B (n_8361), .C (n_8075), .D (n_8588), .Q
       (n_1399));
  NA2X1 g92074(.A (n_7965), .B (n_175), .Q (n_1398));
  AN22X1 g50477(.A (n_8071), .B (n_8361), .C (n_8072), .D (n_8588), .Q
       (n_1397));
  NA2X1 g92075(.A (n_7963), .B (n_175), .Q (n_1396));
  AN22X1 g50468(.A (n_8069), .B (n_8361), .C (n_8070), .D (n_8588), .Q
       (n_1395));
  NA2X1 g92076(.A (n_7962), .B (n_175), .Q (n_1394));
  AN22X1 g50484(.A (n_8067), .B (n_8361), .C (n_8068), .D (n_8588), .Q
       (n_1393));
  NA2X1 g92077(.A (n_7961), .B (n_175), .Q (n_1392));
  AN22X1 g50478(.A (n_8065), .B (n_8361), .C (n_8066), .D (n_8588), .Q
       (n_1391));
  NA2X1 g92078(.A (n_7960), .B (n_175), .Q (n_1390));
  AN22X1 g50469(.A (n_8063), .B (n_8361), .C (n_8064), .D (n_8588), .Q
       (n_1389));
  NA2X1 g92079(.A (n_7959), .B (n_175), .Q (n_1388));
  AN22X1 g50460(.A (n_8061), .B (n_8361), .C (n_8062), .D (n_8588), .Q
       (n_1387));
  NA2X1 g92080(.A (n_7958), .B (n_175), .Q (n_1386));
  AN22X1 g50491(.A (n_8059), .B (n_8361), .C (n_8060), .D (n_8588), .Q
       (n_1385));
  NA2X1 g92081(.A (n_7957), .B (n_175), .Q (n_1384));
  AN22X1 g50487(.A (n_8057), .B (n_8361), .C (n_8058), .D (n_8588), .Q
       (n_1383));
  AN222X1 g50345(.A (n_8149), .B (n_8361), .C (n_8150), .D (n_8588), .E
       (n_8003), .F (n_8587), .Q (n_1382));
  NA2X1 g92082(.A (n_7949), .B (n_175), .Q (n_1381));
  AN22X1 g50474(.A (n_8055), .B (n_8361), .C (n_8056), .D (n_8588), .Q
       (n_1380));
  NA2X1 g92083(.A (n_7928), .B (n_175), .Q (n_1379));
  AN22X1 g50465(.A (n_8050), .B (n_8361), .C (n_8052), .D (n_8588), .Q
       (n_1378));
  NA2X1 g92084(.A (n_7924), .B (n_175), .Q (n_1377));
  AN22X1 g50486(.A (n_8038), .B (n_8361), .C (n_8044), .D (n_8588), .Q
       (n_1376));
  NA2X1 g92085(.A (n_7922), .B (n_175), .Q (n_1375));
  AN22X1 g50475(.A (n_8027), .B (n_8361), .C (n_8032), .D (n_8588), .Q
       (n_1374));
  NA2X1 g92086(.A (n_7921), .B (n_175), .Q (n_1373));
  AN22X1 g50467(.A (n_8025), .B (n_8361), .C (n_8026), .D (n_8588), .Q
       (n_1372));
  AN22X1 g50457(.A (n_8352), .B (n_8361), .C (n_8024), .D (n_8588), .Q
       (n_1370));
  NA2X1 g92088(.A (n_7919), .B (n_175), .Q (n_1369));
  AN22X1 g50476(.A (n_8021), .B (n_8361), .C (n_8022), .D (n_8588), .Q
       (n_1368));
  NA2X1 g92089(.A (n_7918), .B (n_175), .Q (n_1367));
  AN22X1 g50466(.A (n_8019), .B (n_8361), .C (n_8020), .D (n_8588), .Q
       (n_1366));
  NA2X1 g92090(.A (n_7917), .B (n_175), .Q (n_1365));
  AN22X1 g50458(.A (n_8017), .B (n_8361), .C (n_8018), .D (n_8588), .Q
       (n_1364));
  NA2X1 g92091(.A (n_7916), .B (n_175), .Q (n_1363));
  AN22X1 g50451(.A (n_8015), .B (n_8361), .C (n_8016), .D (n_8588), .Q
       (n_1362));
  AN222X1 g50340(.A (n_8147), .B (n_8361), .C (n_8148), .D (n_8588), .E
       (n_8002), .F (n_8587), .Q (n_1361));
  NA2X1 g92092(.A (n_7915), .B (n_175), .Q (n_1360));
  AN22X1 g50452(.A (n_8013), .B (n_8361), .C (n_8014), .D (n_8588), .Q
       (n_1359));
  AN21X1 g50247(.A (n_7914), .B (n_175), .C (n_1102), .Q (n_1358));
  NA2X1 g92093(.A (n_7913), .B (n_175), .Q (n_1357));
  AN22X1 g50443(.A (n_8009), .B (n_8361), .C (n_8010), .D (n_8588), .Q
       (n_1356));
  AN22X1 g50441(.A (n_8351), .B (n_8361), .C (n_8008), .D (n_8588), .Q
       (n_1354));
  AN222X1 g50333(.A (n_8145), .B (n_8361), .C (n_8146), .D (n_8588), .E
       (n_8001), .F (n_8587), .Q (n_1353));
  AN222X1 g50310(.A (n_8143), .B (n_8361), .C (n_8144), .D (n_8588), .E
       (n_8000), .F (n_8587), .Q (n_1352));
  AN222X1 g50311(.A (n_8141), .B (n_8361), .C (n_8142), .D (n_8588), .E
       (n_7999), .F (n_8587), .Q (n_1351));
  AN222X1 g50306(.A (n_8139), .B (n_8361), .C (n_8140), .D (n_8588), .E
       (n_7998), .F (n_8587), .Q (n_1350));
  NA2X1 g92095(.A (n_1169), .B (n_8354), .Q (n_1349));
  NA2X1 g92096(.A (take_trap_39229), .B (program_counter[10]), .Q
       (n_1348));
  NA2X1 g92097(.A (n_1169), .B (n_7395), .Q (n_1347));
  NA2X1 g92098(.A (take_trap_39229), .B (program_counter[11]), .Q
       (n_1346));
  NA2X1 g92099(.A (n_1169), .B (n_7394), .Q (n_1345));
  NA2X1 g92100(.A (take_trap_39229), .B (program_counter[12]), .Q
       (n_1344));
  NA2X1 g92101(.A (n_1169), .B (n_7393), .Q (n_1343));
  NA2X1 g92102(.A (take_trap_39229), .B (program_counter[13]), .Q
       (n_1342));
  NA2X1 g92103(.A (n_1169), .B (n_7392), .Q (n_1341));
  NA2X1 g92104(.A (take_trap_39229), .B (program_counter[14]), .Q
       (n_1340));
  NA2X1 g92105(.A (n_1169), .B (n_7391), .Q (n_1339));
  NA2X1 g92106(.A (take_trap_39229), .B (program_counter[15]), .Q
       (n_1338));
  NA2X1 g92107(.A (n_1169), .B (n_8622), .Q (n_1337));
  NA2X1 g92108(.A (take_trap_39229), .B (program_counter[16]), .Q
       (n_1336));
  NA2X1 g92109(.A (n_1169), .B (n_7389), .Q (n_1335));
  NA2X1 g92110(.A (take_trap_39229), .B (program_counter[17]), .Q
       (n_1334));
  NA2X1 g92111(.A (n_1169), .B (n_7388), .Q (n_1333));
  NA2X1 g92112(.A (take_trap_39229), .B (program_counter[18]), .Q
       (n_1332));
  NA2X1 g92113(.A (n_1169), .B (n_7387), .Q (n_1331));
  NA2X1 g92114(.A (take_trap_39229), .B (program_counter[19]), .Q
       (n_1330));
  NA2X1 g92115(.A (n_1169), .B (n_7386), .Q (n_1329));
  NA2X1 g92116(.A (take_trap_39229), .B (program_counter[20]), .Q
       (n_1328));
  NA2X1 g92117(.A (n_1169), .B (n_7385), .Q (n_1327));
  NA2X1 g92118(.A (take_trap_39229), .B (program_counter[21]), .Q
       (n_1326));
  NA2X1 g92119(.A (n_1169), .B (n_7384), .Q (n_1325));
  NA2X1 g92120(.A (take_trap_39229), .B (program_counter[22]), .Q
       (n_1324));
  NA2X1 g92121(.A (n_1169), .B (n_7383), .Q (n_1323));
  NA2X1 g92122(.A (take_trap_39229), .B (program_counter[23]), .Q
       (n_1322));
  NA2X1 g92123(.A (n_1169), .B (n_8571), .Q (n_1321));
  NA2X1 g92124(.A (take_trap_39229), .B (program_counter[24]), .Q
       (n_1320));
  NA2X1 g92125(.A (n_1169), .B (n_7381), .Q (n_1319));
  NA2X1 g92126(.A (take_trap_39229), .B (program_counter[25]), .Q
       (n_1318));
  NA2X1 g92127(.A (n_1169), .B (n_7380), .Q (n_1317));
  NA2X1 g92128(.A (take_trap_39229), .B (program_counter[26]), .Q
       (n_1316));
  NA2X1 g92129(.A (n_1169), .B (n_7379), .Q (n_1315));
  NA2X1 g92130(.A (take_trap_39229), .B (program_counter[27]), .Q
       (n_1314));
  NA2X1 g92131(.A (n_1169), .B (n_7378), .Q (n_1313));
  NA2X1 g92132(.A (take_trap_39229), .B (program_counter[28]), .Q
       (n_1312));
  NA2X1 g92133(.A (n_1169), .B (n_7377), .Q (n_1311));
  NA2X1 g92134(.A (take_trap_39229), .B (program_counter[29]), .Q
       (n_1310));
  NA2X1 g92135(.A (n_1169), .B (n_6233), .Q (n_1309));
  NA2X1 g92136(.A (take_trap_39229), .B (program_counter[2]), .Q
       (n_1308));
  NA2X1 g92137(.A (n_1169), .B (n_7376), .Q (n_1307));
  NA2X1 g92138(.A (take_trap_39229), .B (program_counter[30]), .Q
       (n_1306));
  NA2X1 g92139(.A (n_1169), .B (n_7635), .Q (n_1305));
  NA2X1 g92140(.A (take_trap_39229), .B (program_counter[31]), .Q
       (n_1304));
  NA2X1 g92141(.A (n_1169), .B (n_6234), .Q (n_1303));
  NA2X1 g92142(.A (take_trap_39229), .B (program_counter[3]), .Q
       (n_1302));
  NA2X1 g92143(.A (n_1169), .B (n_7632), .Q (n_1301));
  NA2X1 g92144(.A (take_trap_39229), .B (program_counter[4]), .Q
       (n_1300));
  NA2X1 g92145(.A (n_1169), .B (n_6232), .Q (n_1299));
  NA2X1 g92146(.A (take_trap_39229), .B (program_counter[5]), .Q
       (n_1298));
  NA2X1 g92147(.A (n_1169), .B (n_6237), .Q (n_1297));
  NA2X1 g92148(.A (take_trap_39229), .B (program_counter[6]), .Q
       (n_1296));
  NA2X1 g92149(.A (n_1169), .B (n_6238), .Q (n_1295));
  NA2X1 g92150(.A (take_trap_39229), .B (program_counter[7]), .Q
       (n_1294));
  NA2X1 g92151(.A (n_1169), .B (n_7398), .Q (n_1293));
  NA2X1 g92152(.A (take_trap_39229), .B (program_counter[8]), .Q
       (n_1292));
  NA2X1 g92153(.A (n_1169), .B (n_7397), .Q (n_1291));
  NA2X1 g92154(.A (take_trap_39229), .B (program_counter[9]), .Q
       (n_1290));
  AN222X1 g50353(.A (n_7592), .B (n_1101), .C (n_7593), .D (n_1100), .E
       (n_7465), .F (n_174), .Q (n_1289));
  AN222X1 g50300(.A (n_7572), .B (n_1101), .C (n_7573), .D (n_1100), .E
       (n_7455), .F (n_174), .Q (n_1288));
  AN222X1 g50296(.A (n_7570), .B (n_1101), .C (n_7571), .D (n_1100), .E
       (n_7454), .F (n_174), .Q (n_1287));
  AN222X1 g50304(.A (n_7568), .B (n_1101), .C (n_7569), .D (n_1100), .E
       (n_7453), .F (n_174), .Q (n_1286));
  AN222X1 g50301(.A (n_7566), .B (n_1101), .C (n_7567), .D (n_1100), .E
       (n_7452), .F (n_174), .Q (n_1285));
  AN222X1 g50297(.A (n_7564), .B (n_1101), .C (n_7565), .D (n_1100), .E
       (n_7451), .F (n_174), .Q (n_1284));
  AN222X1 g50292(.A (n_1101), .B (n_7562), .C (n_7563), .D (n_1100), .E
       (n_159), .F (n_7450), .Q (n_1283));
  AN222X1 g50293(.A (n_1101), .B (n_7560), .C (n_1100), .D (n_7561), .E
       (n_159), .F (n_7449), .Q (n_1282));
  AN222X1 g50286(.A (n_1101), .B (n_7558), .C (n_1100), .D (n_7559), .E
       (n_159), .F (n_7448), .Q (n_1281));
  AN222X1 g50279(.A (n_1101), .B (n_7556), .C (n_1100), .D (n_7557), .E
       (n_159), .F (n_7447), .Q (n_1280));
  AN222X1 g50274(.A (n_7554), .B (n_1101), .C (n_1100), .D (n_7555), .E
       (n_159), .F (n_7446), .Q (n_1279));
  AN222X1 g50350(.A (n_7590), .B (n_1101), .C (n_7591), .D (n_1100), .E
       (n_7464), .F (n_174), .Q (n_1278));
  AN222X1 g50287(.A (n_1101), .B (n_7552), .C (n_1100), .D (n_7553), .E
       (n_159), .F (n_7445), .Q (n_1277));
  AN222X1 g50280(.A (n_1101), .B (n_7550), .C (n_1100), .D (n_7551), .E
       (n_159), .F (n_7444), .Q (n_1276));
  AN222X1 g50288(.A (n_1101), .B (n_7548), .C (n_1100), .D (n_7549), .E
       (n_159), .F (n_7443), .Q (n_1275));
  AN222X1 g50281(.A (n_1101), .B (n_7546), .C (n_1100), .D (n_7547), .E
       (n_159), .F (n_7442), .Q (n_1274));
  AN222X1 g50289(.A (n_1101), .B (n_7544), .C (n_1100), .D (n_7545), .E
       (n_159), .F (n_7441), .Q (n_1273));
  AN222X1 g50282(.A (n_1101), .B (n_7542), .C (n_1100), .D (n_7543), .E
       (n_159), .F (n_7440), .Q (n_1272));
  AN222X1 g50275(.A (n_7540), .B (n_1101), .C (n_1100), .D (n_7541), .E
       (n_159), .F (n_7439), .Q (n_1271));
  AN222X1 g50270(.A (n_7538), .B (n_1101), .C (n_1100), .D (n_7539), .E
       (n_159), .F (n_7438), .Q (n_1270));
  AN222X1 g50271(.A (n_1101), .B (n_7536), .C (n_1100), .D (n_7537), .E
       (n_159), .F (n_7437), .Q (n_1269));
  AN222X1 g50267(.A (n_7534), .B (n_1101), .C (n_1100), .D (n_7535), .E
       (n_159), .F (n_8349), .Q (n_1268));
  AN222X1 g50347(.A (n_7588), .B (n_1101), .C (n_7589), .D (n_1100), .E
       (n_7463), .F (n_174), .Q (n_1267));
  AN21X1 g50265(.A (n_7435), .B (n_159), .C (n_1099), .Q (n_1266));
  AN22X1 g50546(.A (n_7530), .B (n_1101), .C (n_7531), .D (n_1100), .Q
       (n_1264));
  AN21X1 g50262(.A (n_7433), .B (n_159), .C (n_1098), .Q (n_1263));
  AN22X1 g50520(.A (n_7526), .B (n_1101), .C (n_7527), .D (n_1100), .Q
       (n_1261));
  AN21X1 g50257(.A (n_7431), .B (n_159), .C (n_1097), .Q (n_1260));
  AN22X1 g50508(.A (n_7522), .B (n_1101), .C (n_7523), .D (n_1100), .Q
       (n_1258));
  NA2X1 g92158(.A (n_7429), .B (n_159), .Q (n_1257));
  AN22X1 g50518(.A (n_7520), .B (n_1101), .C (n_7521), .D (n_1100), .Q
       (n_1256));
  NA2X1 g92159(.A (n_7427), .B (n_159), .Q (n_1254));
  AN22X1 g50548(.A (n_7516), .B (n_1101), .C (n_7517), .D (n_1100), .Q
       (n_1253));
  AN222X1 g50344(.A (n_7586), .B (n_1101), .C (n_7587), .D (n_1100), .E
       (n_7462), .F (n_174), .Q (n_1251));
  NA2X1 g92160(.A (n_7425), .B (n_159), .Q (n_1250));
  AN22X1 g50510(.A (n_7512), .B (n_1101), .C (n_7513), .D (n_1100), .Q
       (n_1249));
  NA2X1 g92161(.A (n_7423), .B (n_159), .Q (n_1247));
  AN22X1 g50482(.A (n_7508), .B (n_1101), .C (n_7509), .D (n_1100), .Q
       (n_1246));
  NA2X1 g92162(.A (n_7420), .B (n_159), .Q (n_1243));
  AN22X1 g50480(.A (n_7502), .B (n_1101), .C (n_7503), .D (n_1100), .Q
       (n_1242));
  NA2X1 g92163(.A (n_7418), .B (n_159), .Q (n_1240));
  AN22X1 g50462(.A (n_7498), .B (n_1101), .C (n_7499), .D (n_1100), .Q
       (n_1239));
  NA2X1 g92164(.A (n_7416), .B (n_159), .Q (n_1237));
  AN22X1 g50472(.A (n_7494), .B (n_1101), .C (n_7495), .D (n_1100), .Q
       (n_1236));
  AN222X1 g50343(.A (n_7584), .B (n_1101), .C (n_7585), .D (n_1100), .E
       (n_7461), .F (n_174), .Q (n_1235));
  NA2X1 g92165(.A (n_7414), .B (n_159), .Q (n_1233));
  AN22X1 g50453(.A (n_7490), .B (n_1101), .C (n_7491), .D (n_1100), .Q
       (n_1232));
  NA2X1 g92166(.A (n_7413), .B (n_159), .Q (n_1231));
  AN22X1 g50473(.A (n_7488), .B (n_1101), .C (n_7489), .D (n_1100), .Q
       (n_1230));
  AN21X1 g50256(.A (n_7412), .B (n_159), .C (n_1088), .Q (n_1229));
  AN22X1 g50454(.A (n_7484), .B (n_1101), .C (n_7485), .D (n_1100), .Q
       (n_1227));
  NA2X1 g92168(.A (n_7408), .B (n_159), .Q (n_1224));
  AN22X1 g50455(.A (n_7478), .B (n_1101), .C (n_7479), .D (n_1100), .Q
       (n_1223));
  AN21X1 g50249(.A (n_7407), .B (n_159), .C (n_1085), .Q (n_1222));
  NA2X1 g92169(.A (n_7406), .B (n_159), .Q (n_1221));
  AN22X1 g50444(.A (n_7474), .B (n_1101), .C (n_7475), .D (n_1100), .Q
       (n_1220));
  AN222X1 g50337(.A (n_7582), .B (n_1101), .C (n_7583), .D (n_1100), .E
       (n_7460), .F (n_174), .Q (n_1219));
  AN22X1 g50445(.A (n_7472), .B (n_1101), .C (n_8350), .D (n_1100), .Q
       (n_1217));
  AN21X1 g50248(.A (n_7404), .B (n_159), .C (n_1084), .Q (n_1216));
  AN22X1 g50439(.A (n_7468), .B (n_1101), .C (n_7469), .D (n_1100), .Q
       (n_1214));
  AN22X1 g50438(.A (n_8353), .B (n_1101), .C (n_7467), .D (n_1100), .Q
       (n_1212));
  AN222X1 g50314(.A (n_7580), .B (n_1101), .C (n_7581), .D (n_1100), .E
       (n_7459), .F (n_174), .Q (n_1211));
  AN222X1 g50308(.A (n_7578), .B (n_1101), .C (n_7579), .D (n_1100), .E
       (n_7458), .F (n_174), .Q (n_1210));
  AN222X1 g50309(.A (n_7576), .B (n_1101), .C (n_7577), .D (n_1100), .E
       (n_7457), .F (n_174), .Q (n_1209));
  AN222X1 g50305(.A (n_7574), .B (n_1101), .C (n_7575), .D (n_1100), .E
       (n_7456), .F (n_174), .Q (n_1208));
  INX1 g92172(.A (n_6236), .Q (n_1207));
  INX1 g92173(.A (n_6235), .Q (n_1206));
  MU2IX1 g50527(.S (n_8340), .IN0 (n_1083), .IN1 (n_7275), .Q (n_1205));
  AN31X1 g92175(.A (n_7249), .B (n_156), .C (n_1447), .D (n_8340), .Q
       (n_1203));
  AN21X1 g50436(.A (n_158), .B (program_counter[0]), .C (n_1080), .Q
       (n_1202));
  AN211X1 g50606(.A (n_158), .B (program_counter[10]), .C (n_1079), .D
       (n_1078), .Q (n_1201));
  AN211X1 g50607(.A (n_158), .B (program_counter[11]), .C (n_1077), .D
       (n_1076), .Q (n_1200));
  AN211X1 g50608(.A (n_158), .B (program_counter[12]), .C (n_1075), .D
       (n_1074), .Q (n_1199));
  AN211X1 g50609(.A (n_158), .B (program_counter[13]), .C (n_1073), .D
       (n_1072), .Q (n_1198));
  AN211X1 g50601(.A (n_158), .B (program_counter[14]), .C (n_1071), .D
       (n_1070), .Q (n_1197));
  AN211X1 g50610(.A (n_158), .B (program_counter[15]), .C (n_1069), .D
       (n_1068), .Q (n_1196));
  AN211X1 g50604(.A (n_158), .B (program_counter[16]), .C (n_1067), .D
       (n_1066), .Q (n_1195));
  AN211X1 g50611(.A (n_158), .B (program_counter[17]), .C (n_1065), .D
       (n_1064), .Q (n_1194));
  AN211X1 g50626(.A (n_158), .B (program_counter[18]), .C (n_1063), .D
       (n_1062), .Q (n_1193));
  AN211X1 g50620(.A (n_158), .B (program_counter[19]), .C (n_1061), .D
       (n_1060), .Q (n_1192));
  AN21X1 g50435(.A (n_158), .B (program_counter[1]), .C (n_1059), .Q
       (n_1191));
  AN211X1 g50612(.A (n_158), .B (program_counter[20]), .C (n_1058), .D
       (n_1057), .Q (n_1190));
  AN211X1 g50613(.A (n_158), .B (program_counter[21]), .C (n_1056), .D
       (n_1055), .Q (n_1189));
  AN211X1 g50614(.A (n_158), .B (program_counter[22]), .C (n_1054), .D
       (n_1053), .Q (n_1188));
  AN211X1 g50615(.A (n_158), .B (program_counter[23]), .C (n_1052), .D
       (n_1051), .Q (n_1187));
  AN211X1 g50605(.A (n_158), .B (program_counter[24]), .C (n_1050), .D
       (n_1049), .Q (n_1186));
  AN211X1 g50616(.A (n_158), .B (program_counter[25]), .C (n_1048), .D
       (n_1047), .Q (n_1185));
  AN211X1 g50617(.A (n_158), .B (program_counter[26]), .C (n_1046), .D
       (n_1045), .Q (n_1184));
  AN211X1 g50602(.A (n_158), .B (program_counter[27]), .C (n_1044), .D
       (n_1043), .Q (n_1183));
  AN211X1 g50618(.A (n_158), .B (program_counter[28]), .C (n_1042), .D
       (n_1041), .Q (n_1182));
  AN211X1 g50603(.A (n_158), .B (program_counter[29]), .C (n_1040), .D
       (n_1039), .Q (n_1181));
  AN211X1 g50599(.A (n_158), .B (program_counter[2]), .C (n_1038), .D
       (n_1037), .Q (n_1180));
  AN211X1 g50600(.A (n_158), .B (program_counter[30]), .C (n_1036), .D
       (n_1035), .Q (n_1179));
  AN211X1 g50619(.A (n_158), .B (program_counter[31]), .C (n_1034), .D
       (n_1033), .Q (n_1178));
  AN211X1 g50621(.A (n_158), .B (program_counter[3]), .C (n_1032), .D
       (n_1031), .Q (n_1177));
  AN211X1 g50622(.A (n_158), .B (program_counter[4]), .C (n_1030), .D
       (n_1029), .Q (n_1176));
  AN211X1 g50598(.A (n_158), .B (program_counter[5]), .C (n_1028), .D
       (n_1027), .Q (n_1175));
  AN211X1 g50623(.A (n_158), .B (program_counter[6]), .C (n_1026), .D
       (n_1025), .Q (n_1174));
  AN211X1 g50624(.A (n_158), .B (program_counter[7]), .C (n_1024), .D
       (n_1023), .Q (n_1173));
  AN211X1 g50625(.A (n_158), .B (program_counter[8]), .C (n_1022), .D
       (n_1021), .Q (n_1172));
  AN211X1 g50597(.A (n_158), .B (program_counter[9]), .C (n_1020), .D
       (n_1019), .Q (n_1171));
  AN21X1 g92176(.A (n_1169), .B (n_1018), .C (flush_37557), .Q
       (n_1170));
  INX4 g51952(.A (take_trap_39229), .Q (n_1169));
  AN221X4 g48169(.A (program_counter[0]), .B (n_2548), .C (n_1017), .D
       (n_155), .E (n_1016), .Q (n_1167));
  AN221X1 g48171(.A (n_1015), .B (n_1014), .C (n_1013), .D (n_7721), .E
       (n_1012), .Q (n_1166));
  AND3X2 g48831(.A (n_1011), .B (n_1010), .C (n_1009), .Q (n_1165));
  AN21X4 g48832(.A (n_7719), .B (n_1013), .C (n_1008), .Q (n_1164));
  AN21X4 g49696(.A (n_7718), .B (n_1013), .C (n_1007), .Q (n_1163));
  AN21X1 g49489(.A (n_7717), .B (n_1013), .C (n_1006), .Q (n_1162));
  AN21X1 g48170(.A (n_7716), .B (n_1013), .C (n_1005), .Q (n_1161));
  AND2X1 g48830(.A (n_1004), .B (n_1003), .Q (n_1160));
  INX3 g49594(.A (n_1002), .Q (n_1159));
  INX4 g49593(.A (n_1001), .Q (n_1158));
  INX4 g49596(.A (n_1000), .Q (n_1157));
  OA211X1 g49488(.A (n_999), .B (n_998), .C (n_997), .D (n_996), .Q
       (n_1156));
  INX3 g48657(.A (n_995), .Q (n_1155));
  INX4 g49595(.A (n_994), .Q (n_1154));
  INX4 g48658(.A (n_993), .Q (n_1153));
  INX4 g49705(.A (n_991), .Q (n_1151));
  INX4 g49708(.A (n_990), .Q (n_1150));
  INX4 g49707(.A (n_989), .Q (n_1149));
  INX4 g49706(.A (n_988), .Q (n_1148));
  INX6 g49597(.A (n_987), .Q (n_1147));
  INX4 g49709(.A (n_986), .Q (n_1146));
  OA211X1 g48829(.A (n_985), .B (n_998), .C (n_984), .D (n_983), .Q
       (n_1145));
  INX6 g49599(.A (n_982), .Q (n_1144));
  INX4 g49598(.A (n_981), .Q (n_1143));
  OA211X1 g49703(.A (n_980), .B (n_998), .C (n_979), .D (n_978), .Q
       (n_1142));
  OA211X1 g48828(.A (n_977), .B (n_998), .C (n_976), .D (n_975), .Q
       (n_1141));
  AND3X2 g48167(.A (n_974), .B (n_973), .C (n_972), .Q (n_1140));
  AND3X1 g48168(.A (n_971), .B (n_970), .C (n_969), .Q (n_1139));
  AN221X1 g48166(.A (n_968), .B (n_967), .C (n_1013), .D (n_7724), .E
       (n_966), .Q (n_1138));
  AN21X1 g48835(.A (n_7723), .B (n_1013), .C (n_965), .Q (n_1137));
  AND3X1 g48833(.A (n_964), .B (n_963), .C (n_962), .Q (n_1136));
  INX1 g92178(.A (n_7609), .Q (n_1135));
  INX1 g92179(.A (n_7608), .Q (n_1134));
  INX1 g92180(.A (n_7607), .Q (n_1133));
  INX1 g92181(.A (n_7605), .Q (n_1132));
  INX1 g92182(.A (n_7604), .Q (n_1131));
  INX1 g92183(.A (n_7603), .Q (n_1130));
  INX1 g92184(.A (n_7602), .Q (n_1129));
  INX1 g92185(.A (n_7601), .Q (n_1128));
  INX1 g92186(.A (n_7600), .Q (n_1127));
  INX1 g92187(.A (n_7599), .Q (n_1126));
  INX1 g92188(.A (n_7598), .Q (n_1125));
  INX1 g92189(.A (n_7597), .Q (n_1124));
  INX1 g92190(.A (n_7596), .Q (n_1123));
  INX1 g92191(.A (n_7624), .Q (n_1122));
  INX1 g92192(.A (n_7623), .Q (n_1121));
  INX1 g92193(.A (n_7622), .Q (n_1120));
  INX1 g92194(.A (n_7621), .Q (n_1119));
  INX1 g92195(.A (n_7620), .Q (n_1118));
  INX1 g92196(.A (n_7619), .Q (n_1117));
  INX1 g92197(.A (n_7617), .Q (n_1116));
  INX1 g92198(.A (n_7618), .Q (n_1115));
  INX1 g92199(.A (n_7606), .Q (n_1114));
  INX1 g92200(.A (n_7627), .Q (n_1113));
  INX1 g92201(.A (n_7616), .Q (n_1112));
  INX1 g92202(.A (n_7615), .Q (n_1111));
  INX1 g92203(.A (n_7614), .Q (n_1110));
  INX1 g92204(.A (n_7613), .Q (n_1109));
  INX1 g92205(.A (n_7612), .Q (n_1108));
  INX1 g92206(.A (n_7611), .Q (n_1107));
  INX1 g92207(.A (n_7610), .Q (n_1106));
  INX6 g52018(.A (n_181), .Q (n_179));
  NO2X1 g92208(.A (n_8361), .B (n_8588), .Q (n_1105));
  BUCX6 g92211(.A (n_8587), .Q (n_175));
  AO22X1 g50448(.A (n_8011), .B (n_8361), .C (n_8012), .D (n_8588), .Q
       (n_1102));
  ON21X4 g92212(.A (n_174), .B (n_7694), .C (n_8157), .Q (n_1101));
  AND2X4 g92213(.A (n_8157), .B (n_7694), .Q (n_1100));
  AO22X1 g50559(.A (n_7532), .B (n_1101), .C (n_7533), .D (n_1100), .Q
       (n_1099));
  BUCX6 g92214(.A (n_174), .Q (n_159));
  AO22X1 g50533(.A (n_7528), .B (n_1101), .C (n_7529), .D (n_1100), .Q
       (n_1098));
  AO22X1 g50513(.A (n_7524), .B (n_1101), .C (n_7525), .D (n_1100), .Q
       (n_1097));
  AO22X1 g50463(.A (n_7486), .B (n_1101), .C (n_7487), .D (n_1100), .Q
       (n_1088));
  AO22X1 g50450(.A (n_7476), .B (n_1101), .C (n_7477), .D (n_1100), .Q
       (n_1085));
  AO22X1 g50442(.A (n_7470), .B (n_1101), .C (n_7471), .D (n_1100), .Q
       (n_1084));
  AO21X1 g92215(.A (n_6256), .B (n_960), .C (n_6234), .Q (n_1083));
  NO2X1 g92216(.A (n_959), .B (n_7714), .Q (n_1082));
  AN21X1 g92217(.A (n_8078), .B (n_7249), .C (n_7714), .Q (n_1081));
  ON22X1 g50627(.A (n_8666), .B (n_958), .C (take_trap_39229), .D
       (n_1207), .Q (n_1080));
  INX1 g92218(.A (n_1349), .Q (n_1079));
  NO2I1X1 g92219(.B (n_8666), .AN (n_7270), .Q (n_1078));
  INX1 g92220(.A (n_1347), .Q (n_1077));
  NO2I1X1 g92221(.B (n_8666), .AN (n_7274), .Q (n_1076));
  INX1 g92222(.A (n_1345), .Q (n_1075));
  NO2I1X1 g92223(.B (n_8666), .AN (n_7277), .Q (n_1074));
  INX1 g92224(.A (n_1343), .Q (n_1073));
  NO2I1X1 g92225(.B (n_8666), .AN (n_7269), .Q (n_1072));
  INX1 g92226(.A (n_1341), .Q (n_1071));
  NO2I1X1 g92227(.B (n_8666), .AN (n_7268), .Q (n_1070));
  INX1 g92228(.A (n_1339), .Q (n_1069));
  NO2I1X1 g92229(.B (n_8666), .AN (n_7267), .Q (n_1068));
  INX1 g92230(.A (n_1337), .Q (n_1067));
  NO2I1X1 g92231(.B (n_8666), .AN (n_7265), .Q (n_1066));
  INX1 g92232(.A (n_1335), .Q (n_1065));
  NO2I1X1 g92233(.B (n_8666), .AN (n_7264), .Q (n_1064));
  INX1 g92234(.A (n_1333), .Q (n_1063));
  NO2I1X1 g92235(.B (n_8666), .AN (n_7263), .Q (n_1062));
  INX1 g92236(.A (n_1331), .Q (n_1061));
  NO2I1X1 g92237(.B (n_8666), .AN (n_7262), .Q (n_1060));
  ON22X1 g50628(.A (n_8666), .B (n_957), .C (take_trap_39229), .D
       (n_1206), .Q (n_1059));
  INX1 g92238(.A (n_1329), .Q (n_1058));
  NO2I1X1 g92239(.B (n_8666), .AN (n_7261), .Q (n_1057));
  INX1 g92240(.A (n_1327), .Q (n_1056));
  NO2I1X1 g92241(.B (n_8666), .AN (n_7260), .Q (n_1055));
  INX1 g92242(.A (n_1325), .Q (n_1054));
  NO2I1X1 g92243(.B (n_8666), .AN (n_7259), .Q (n_1053));
  INX1 g92244(.A (n_1323), .Q (n_1052));
  NO2I1X1 g92245(.B (n_8666), .AN (n_7258), .Q (n_1051));
  INX1 g92246(.A (n_1321), .Q (n_1050));
  NO2I1X1 g92247(.B (n_8666), .AN (n_7257), .Q (n_1049));
  INX1 g92248(.A (n_1319), .Q (n_1048));
  NO2I1X1 g92249(.B (n_8666), .AN (n_7256), .Q (n_1047));
  INX1 g92250(.A (n_1317), .Q (n_1046));
  NO2I1X1 g92251(.B (n_8666), .AN (n_7255), .Q (n_1045));
  INX1 g92252(.A (n_1315), .Q (n_1044));
  NO2I1X1 g92253(.B (n_8666), .AN (n_7254), .Q (n_1043));
  INX1 g92254(.A (n_1313), .Q (n_1042));
  NO2I1X1 g92255(.B (n_8666), .AN (n_7253), .Q (n_1041));
  INX1 g92256(.A (n_1311), .Q (n_1040));
  NO2I1X1 g92257(.B (n_8666), .AN (n_7252), .Q (n_1039));
  INX1 g92258(.A (n_1309), .Q (n_1038));
  NO2I1X1 g92259(.B (n_8666), .AN (n_7280), .Q (n_1037));
  INX1 g92260(.A (n_1307), .Q (n_1036));
  NO2I1X1 g92261(.B (n_8666), .AN (n_7250), .Q (n_1035));
  INX1 g92262(.A (n_1305), .Q (n_1034));
  NO2I1X1 g92263(.B (n_8666), .AN (n_7251), .Q (n_1033));
  INX1 g92264(.A (n_1303), .Q (n_1032));
  NO2I1X1 g92265(.B (n_8666), .AN (n_7279), .Q (n_1031));
  INX1 g92266(.A (n_1301), .Q (n_1030));
  NO2I1X1 g92267(.B (n_8666), .AN (n_7278), .Q (n_1029));
  INX1 g92268(.A (n_1299), .Q (n_1028));
  NO2I1X1 g92269(.B (n_8666), .AN (n_7273), .Q (n_1027));
  INX1 g92270(.A (n_1297), .Q (n_1026));
  NO2I1X1 g92271(.B (n_8666), .AN (n_7272), .Q (n_1025));
  INX1 g92272(.A (n_1295), .Q (n_1024));
  NO2I1X1 g92273(.B (n_8666), .AN (n_7276), .Q (n_1023));
  INX1 g92274(.A (n_1293), .Q (n_1022));
  NO2I1X1 g92275(.B (n_8666), .AN (n_7266), .Q (n_1021));
  INX1 g92276(.A (n_1291), .Q (n_1020));
  NO2I1X1 g92277(.B (n_8666), .AN (n_7271), .Q (n_1019));
  INX1 g92278(.A (n_8523), .Q (n_1018));
  AN211X0 g49816(.A (n_956), .B (n_8309), .C (n_955), .D (n_954), .Q
       (n_1017));
  ON211X1 g49745(.A (n_951), .B (n_998), .C (n_950), .D (n_949), .Q
       (n_1016));
  INX1 g50501(.A (n_948), .Q (n_1015));
  ON22X1 g49959(.A (n_947), .B (alu_2nd_operand[3]), .C (n_946), .D
       (n_945), .Q (n_1014));
  AND2X4 g92279(.A (n_944), .B (n_8163), .Q (n_1013));
  ON211X1 g48722(.A (n_943), .B (n_942), .C (n_941), .D (n_940), .Q
       (n_1012));
  NA2X1 g50446(.A (n_7720), .B (n_1013), .Q (n_1011));
  AN221X1 g49759(.A (n_939), .B (n_938), .C (n_1015), .D (n_937), .E
       (n_154), .Q (n_1010));
  AN221X1 g49688(.A (n_8296), .B (n_7274), .C (n_936), .D (n_935), .E
       (n_934), .Q (n_1009));
  ON211X1 g49299(.A (n_933), .B (n_948), .C (n_932), .D (n_931), .Q
       (n_1008));
  NA3X1 g49723(.A (n_930), .B (n_929), .C (n_928), .Q (n_1007));
  ON211X1 g49694(.A (n_927), .B (n_948), .C (n_926), .D (n_925), .Q
       (n_1006));
  ON21X1 g48594(.A (n_924), .B (n_948), .C (n_923), .Q (n_1005));
  NA2X1 g50440(.A (n_7715), .B (n_1013), .Q (n_1004));
  AN221X1 g49297(.A (n_8296), .B (n_7265), .C (n_922), .D (n_921), .E
       (n_920), .Q (n_1003));
  AO21X2 g49697(.A (n_7713), .B (n_1013), .C (n_919), .Q (n_1002));
  AO21X2 g49695(.A (n_7712), .B (n_1013), .C (n_918), .Q (n_1001));
  AO21X2 g49699(.A (n_7711), .B (n_1013), .C (n_917), .Q (n_1000));
  MU2IX1 g49960(.S (alu_2nd_operand[3]), .IN0 (n_916), .IN1 (n_915), .Q
       (n_999));
  NA2X1 g50589(.A (n_8677), .B (n_914), .Q (n_998));
  AN21X1 g49843(.A (n_913), .B (n_914), .C (n_912), .Q (n_997));
  AN221X1 g49731(.A (read_data[1]), .B (n_911), .C (n_1013), .D
       (n_7730), .E (n_910), .Q (n_996));
  AO21X2 g48834(.A (n_7709), .B (n_1013), .C (n_909), .Q (n_995));
  AO21X2 g49698(.A (n_7706), .B (n_1013), .C (n_908), .Q (n_994));
  AO21X2 g48836(.A (n_7705), .B (n_1013), .C (n_907), .Q (n_993));
  AO21X2 g49717(.A (n_7703), .B (n_1013), .C (n_904), .Q (n_991));
  AO21X2 g49720(.A (n_7702), .B (n_1013), .C (n_903), .Q (n_990));
  AO21X4 g49719(.A (n_7701), .B (n_1013), .C (n_902), .Q (n_989));
  AO21X4 g49718(.A (n_7700), .B (n_1013), .C (n_901), .Q (n_988));
  AO21X2 g49700(.A (n_7699), .B (n_1013), .C (n_900), .Q (n_987));
  AO21X4 g49721(.A (n_7698), .B (n_1013), .C (n_899), .Q (n_986));
  OA222X1 g49955(.A (n_898), .B (n_897), .C (n_896), .D (n_895), .E
       (n_943), .F (n_173), .Q (n_985));
  AN221X1 g49687(.A (n_1013), .B (n_7729), .C (n_894), .D (n_893), .E
       (n_892), .Q (n_984));
  AN211X1 g49847(.A (n_911), .B (read_data[2]), .C (n_891), .D (n_890),
       .Q (n_983));
  AO21X2 g49702(.A (n_7697), .B (n_1013), .C (n_889), .Q (n_982));
  AO21X4 g49701(.A (n_7696), .B (n_1013), .C (n_888), .Q (n_981));
  AN21X1 g49958(.A (n_938), .B (alu_2nd_operand[3]), .C (n_887), .Q
       (n_980));
  AN21X1 g49724(.A (n_7728), .B (n_1013), .C (n_886), .Q (n_979));
  AN21X1 g49840(.A (n_935), .B (n_894), .C (n_885), .Q (n_978));
  AN21X1 g49946(.A (n_884), .B (n_173), .C (n_883), .Q (n_977));
  AN221X1 g49302(.A (n_882), .B (n_881), .C (n_1013), .D (n_7727), .E
       (n_880), .Q (n_976));
  OA221X1 g49894(.A (n_153), .B (n_879), .C (n_878), .D (n_877), .E
       (n_876), .Q (n_975));
  AN21X1 g49803(.A (n_875), .B (n_968), .C (n_874), .Q (n_974));
  NA2X1 g50459(.A (n_7726), .B (n_1013), .Q (n_973));
  AN221X1 g48726(.A (read_data[5]), .B (n_911), .C (n_882), .D (n_873),
       .E (n_872), .Q (n_972));
  AN21X1 g49799(.A (n_871), .B (n_968), .C (n_870), .Q (n_971));
  NA2X1 g50456(.A (n_7725), .B (n_1013), .Q (n_970));
  AN221X1 g48725(.A (read_data[6]), .B (n_911), .C (n_882), .D (n_869),
       .E (n_868), .Q (n_969));
  INX1 g50502(.A (n_998), .Q (n_968));
  ON222X1 g50237(.A (n_898), .B (n_867), .C (n_896), .D (n_866), .E
       (n_865), .F (n_864), .Q (n_967));
  ON211X1 g48723(.A (n_863), .B (n_862), .C (n_861), .D (n_860), .Q
       (n_966));
  ON211X1 g49298(.A (n_859), .B (n_948), .C (n_858), .D (n_857), .Q
       (n_965));
  NA2X1 g50447(.A (n_7722), .B (n_1013), .Q (n_964));
  AN221X1 g49691(.A (n_939), .B (n_915), .C (n_1015), .D (n_856), .E
       (n_855), .Q (n_963));
  AN221X1 g49758(.A (n_8296), .B (n_7271), .C (n_894), .D (n_916), .E
       (n_854), .Q (n_962));
  INX3 g92280(.A (reset_internal_39074), .Q (n_181));
  INX1 g92281(.A (n_8587), .Q (n_178));
  NO2X1 g92284(.A (n_959), .B (n_3869_BAR), .Q (n_174));
  INX1 g51950(.A (n_8157), .Q (n_959));
  NA2I1X1 g92288(.B (n_853), .AN (n_8301), .Q (n_956));
  OR4X1 g92289(.A (n_2548), .B (n_8157), .C (n_4696), .D (n_852), .Q
       (n_955));
  ON221X1 g49846(.A (n_851), .B (n_850), .C (n_849), .D (n_848), .E
       (n_847), .Q (n_954));
  NA2X1 g49301(.A (n_846), .B (n_845), .Q (n_953));
  NO3I1X1 g92290(.B (n_844), .C (n_843), .AN (n_842), .Q (n_952));
  MU2IX1 g49851(.S (alu_2nd_operand[3]), .IN0 (n_841), .IN1 (n_840), .Q
       (n_951));
  AN221X1 g49899(.A (n_839), .B (n_838), .C (n_837), .D (n_836), .E
       (n_835), .Q (n_950));
  AN221X1 g49791(.A (n_834), .B (n_833), .C (read_data[0]), .D (n_911),
       .E (n_832), .Q (n_949));
  NA2X1 g50588(.A (n_831), .B (n_830), .Q (n_948));
  INX1 g50325(.A (n_829), .Q (n_947));
  OA221X2 g92291(.A (n_828), .B (n_827), .C (n_826), .D (n_166), .E
       (n_152), .Q (n_946));
  NA2X1 g92292(.A (n_8496), .B (alu_2nd_operand[3]), .Q (n_945));
  INX1 g92293(.A (n_955), .Q (n_944));
  OA22X1 g50402(.A (n_825), .B (alu_2nd_operand[2]), .C (n_824), .D
       (n_823), .Q (n_943));
  INX1 g50497(.A (n_939), .Q (n_942));
  AN221X1 g49303(.A (n_8296), .B (n_7270), .C (n_936), .D (n_893), .E
       (n_822), .Q (n_941));
  AN21X1 g49832(.A (n_821), .B (alu_2nd_operand[1]), .C (n_820), .Q
       (n_940));
  AND2X1 g50579(.A (n_819), .B (n_914), .Q (n_939));
  ON22X1 g50403(.A (n_866), .B (alu_2nd_operand[2]), .C (n_823), .D
       (n_864), .Q (n_938));
  ON22X1 g49954(.A (n_818), .B (alu_2nd_operand[3]), .C (n_817), .D
       (n_945), .Q (n_937));
  AND2X1 g50585(.A (n_816), .B (n_914), .Q (n_936));
  MU2IX1 g50395(.S (alu_2nd_operand[2]), .IN0 (n_815), .IN1 (n_814), .Q
       (n_935));
  ON221X1 g49751(.A (n_878), .B (n_867), .C (n_813), .D (n_812), .E
       (n_811), .Q (n_934));
  AN21X1 g49957(.A (n_881), .B (alu_2nd_operand[3]), .C (n_810), .Q
       (n_933));
  AN211X1 g49689(.A (n_884), .B (n_894), .C (n_154), .D (n_809), .Q
       (n_932));
  NA2X1 g92294(.A (n_7277), .B (n_8296), .Q (n_931));
  AN221X1 g49806(.A (n_894), .B (n_808), .C (n_1015), .D (n_807), .E
       (n_806), .Q (n_930));
  NA2X1 g92295(.A (n_7269), .B (n_8296), .Q (n_929));
  AN211X1 g49763(.A (n_805), .B (read_data[13]), .C (n_804), .D
       (n_803), .Q (n_928));
  INX1 g49877(.A (n_802), .Q (n_927));
  AN21X1 g49838(.A (n_801), .B (n_894), .C (n_800), .Q (n_926));
  AN211X1 g49727(.A (n_7268), .B (n_8296), .C (n_799), .D (n_803), .Q
       (n_925));
  MU2IX1 g49852(.S (alu_2nd_operand[3]), .IN0 (n_798), .IN1 (n_797), .Q
       (n_924));
  AN221X1 g48724(.A (n_8296), .B (n_7267), .C (n_936), .D (n_796), .E
       (n_795), .Q (n_923));
  INX1 g50504(.A (n_794), .Q (n_922));
  INX1 g49833(.A (n_951), .Q (n_921));
  ON211X1 g49726(.A (n_793), .B (n_792), .C (n_791), .D (n_790), .Q
       (n_920));
  ON211X1 g49713(.A (n_999), .B (n_794), .C (n_789), .D (n_788), .Q
       (n_919));
  NA2X1 g49715(.A (n_787), .B (n_171), .Q (n_918));
  NA2X1 g49711(.A (n_786), .B (n_785), .Q (n_917));
  MU2IX1 g50320(.S (alu_2nd_operand[2]), .IN0 (n_784), .IN1 (n_783), .Q
       (n_916));
  MU2IX1 g50398(.S (alu_2nd_operand[2]), .IN0 (n_782), .IN1 (n_781), .Q
       (n_915));
  NO2X1 g92296(.A (n_955), .B (n_6195), .Q (n_914));
  ON22X1 g50517(.A (n_780), .B (n_779), .C (n_778), .D (n_826), .Q
       (n_913));
  ON321X1 g49900(.A (alu_2nd_operand[0]), .B (n_777), .C (n_776), .D
       (n_878), .E (n_775), .F (n_774), .Q (n_912));
  AO21X1 g92297(.A (n_8165), .B (n_773), .C (n_805), .Q (n_911));
  NA2X1 g49753(.A (n_772), .B (n_771), .Q (n_910));
  AO21X1 g49295(.A (n_7261), .B (n_8296), .C (n_770), .Q (n_909));
  NA2X1 g49728(.A (n_769), .B (n_768), .Q (n_908));
  AO21X1 g49296(.A (n_7259), .B (n_8296), .C (n_767), .Q (n_907));
  NA2X2 g50437(.A (n_7704), .B (n_1013), .Q (n_906));
  AN21X1 g49739(.A (n_7258), .B (n_8296), .C (n_766), .Q (n_905));
  NA3X1 g49735(.A (n_765), .B (n_764), .C (n_763), .Q (n_904));
  NA3X1 g49736(.A (n_762), .B (n_761), .C (n_760), .Q (n_903));
  NA3X1 g49740(.A (n_759), .B (n_758), .C (n_757), .Q (n_902));
  NA3X1 g49738(.A (n_756), .B (n_755), .C (n_754), .Q (n_901));
  NA2X1 g49712(.A (n_753), .B (n_752), .Q (n_900));
  ON211X1 g49737(.A (n_751), .B (n_170), .C (n_750), .D (n_8589), .Q
       (n_899));
  NA2X1 g92298(.A (n_8496), .B (n_173), .Q (n_898));
  AND4X1 g50667(.A (n_748), .B (n_747), .C (n_746), .D (n_745), .Q
       (n_897));
  NA2X1 g92299(.A (alu_2nd_operand[2]), .B (n_173), .Q (n_896));
  AND4X1 g50652(.A (n_744), .B (n_743), .C (n_742), .D (n_741), .Q
       (n_895));
  AND2X1 g50586(.A (n_740), .B (n_914), .Q (n_894));
  MU2X1 g50393(.S (alu_2nd_operand[2]), .IN0 (n_739), .IN1 (n_738), .Q
       (n_893));
  NA3X1 g49754(.A (n_737), .B (n_736), .C (n_735), .Q (n_892));
  ON22X1 g50189(.A (n_946), .B (n_734), .C (n_733), .D (n_732), .Q
       (n_891));
  ON22X1 g50185(.A (n_731), .B (n_153), .C (n_730), .D (n_729), .Q
       (n_890));
  NA2X1 g49710(.A (n_728), .B (n_727), .Q (n_889));
  ON221X1 g49714(.A (n_170), .B (n_726), .C (n_725), .D (n_924), .E
       (n_724), .Q (n_888));
  ON22X1 g50312(.A (n_812), .B (n_898), .C (n_867), .D (n_896), .Q
       (n_887));
  ON211X1 g49746(.A (n_817), .B (n_734), .C (n_723), .D (n_722), .Q
       (n_886));
  ON222X1 g49908(.A (n_721), .B (n_730), .C (n_153), .D (n_720), .E
       (n_733), .F (n_779), .Q (n_885));
  MU2IX1 g50319(.S (alu_2nd_operand[2]), .IN0 (n_719), .IN1 (n_718), .Q
       (n_884));
  NO2X1 g50339(.A (n_717), .B (n_945), .Q (n_883));
  AND2X1 g50584(.A (n_816), .B (n_830), .Q (n_882));
  ON22X1 g50401(.A (n_169), .B (alu_2nd_operand[2]), .C (n_823), .D
       (n_827), .Q (n_881));
  NA3X1 g49732(.A (n_716), .B (n_715), .C (n_714), .Q (n_880));
  AND4X1 g50647(.A (n_713), .B (n_712), .C (n_711), .D (n_710), .Q
       (n_879));
  OR2X1 g50587(.A (n_709), .B (n_708), .Q (n_878));
  AND4X1 g50648(.A (n_707), .B (n_706), .C (n_705), .D (n_704), .Q
       (n_877));
  AN21X1 g50176(.A (n_836), .B (n_703), .C (n_702), .Q (n_876));
  ON22X1 g49952(.A (n_701), .B (alu_2nd_operand[3]), .C (n_781), .D
       (n_945), .Q (n_875));
  ON221X1 g49898(.A (n_153), .B (n_700), .C (n_878), .D (n_784), .E
       (n_699), .Q (n_874));
  ON22X1 g50399(.A (n_168), .B (alu_2nd_operand[2]), .C (n_823), .D
       (n_698), .Q (n_873));
  AO221X1 g49683(.A (n_8296), .B (n_7273), .C (n_697), .D
       (read_data[21]), .E (n_696), .Q (n_872));
  ON22X1 g49948(.A (n_695), .B (alu_2nd_operand[3]), .C (n_865), .D
       (n_824), .Q (n_871));
  ON221X1 g49895(.A (n_776), .B (n_731), .C (n_878), .D (n_897), .E
       (n_694), .Q (n_870));
  MU2IX1 g50400(.S (alu_2nd_operand[2]), .IN0 (n_693), .IN1 (n_946), .Q
       (n_869));
  AO221X1 g49684(.A (n_8296), .B (n_7272), .C (n_697), .D
       (read_data[22]), .E (n_692), .Q (n_868));
  AND4X1 g50668(.A (n_691), .B (n_690), .C (n_689), .D (n_688), .Q
       (n_867));
  OA211X1 g50656(.A (n_687), .B (n_686), .C (n_685), .D (n_684), .Q
       (n_866));
  NA2X1 g92300(.A (n_167), .B (alu_2nd_operand[3]), .Q (n_865));
  NA2X1 g92301(.A (n_683), .B (n_6134), .Q (n_864));
  INX1 g50145(.A (n_797), .Q (n_863));
  INX1 g50500(.A (n_882), .Q (n_862));
  AN21X1 g49884(.A (n_796), .B (n_894), .C (n_682), .Q (n_861));
  AN221X1 g49685(.A (n_773), .B (n_8623), .C (n_8296), .D (n_7276), .E
       (n_680), .Q (n_860));
  OA22X1 g49951(.A (n_793), .B (alu_2nd_operand[3]), .C (n_865), .D
       (n_827), .Q (n_859));
  AN221X1 g49836(.A (n_894), .B (n_841), .C (n_939), .D (n_840), .E
       (n_679), .Q (n_858));
  AN211X1 g49730(.A (n_7266), .B (n_8296), .C (n_678), .D (n_820), .Q
       (n_857));
  ON22X1 g49956(.A (n_677), .B (alu_2nd_operand[3]), .C (n_865), .D
       (n_698), .Q (n_856));
  ON221X1 g49750(.A (n_153), .B (n_775), .C (n_776), .D (n_700), .E
       (n_676), .Q (n_855));
  INX1 g49815(.A (n_940), .Q (n_854));
  AND2X1 g92303(.A (n_674), .B (n_673), .Q (n_853));
  INX1 g92304(.A (n_8073), .Q (n_852));
  AN22X1 g50535(.A (n_672), .B (n_842), .C (n_671), .D (n_670), .Q
       (n_851));
  NA3X1 g50567(.A (n_669), .B (n_668), .C (n_667), .Q (n_850));
  NA2X1 g92305(.A (n_666), .B (n_665), .Q (n_849));
  AN22X1 g50536(.A (n_664), .B (n_663), .C (n_662), .D (n_661), .Q
       (n_848));
  AN222X1 g50191(.A (n_666), .B (n_660), .C (n_673), .D (n_659), .E
       (n_658), .F (n_669), .Q (n_847));
  NA3X1 g49690(.A (n_657), .B (n_656), .C (n_655), .Q (n_846));
  AN22X1 g50540(.A (n_656), .B (n_654), .C (n_653), .D (n_652), .Q
       (n_845));
  NO2I1X1 g92306(.B (n_6132), .AN (n_8495), .Q (n_844));
  AND2X1 g92307(.A (alu_2nd_operand[17]), .B (n_651), .Q (n_843));
  AN21X1 g92308(.A (alu_2nd_operand[18]), .B (n_650), .C (n_649), .Q
       (n_842));
  MU2IX1 g50316(.S (alu_2nd_operand[2]), .IN0 (n_877), .IN1 (n_719), .Q
       (n_841));
  MU2IX1 g50240(.S (alu_2nd_operand[2]), .IN0 (n_718), .IN1 (n_717), .Q
       (n_840));
  NO2X1 g50590(.A (n_648), .B (n_708), .Q (n_839));
  INX1 g50595(.A (n_879), .Q (n_838));
  INX1 g50506(.A (n_153), .Q (n_837));
  ON211X1 g50571(.A (n_729), .B (alu_2nd_operand[1]), .C (n_647), .D
       (n_646), .Q (n_836));
  ON22X1 g50180(.A (n_645), .B (n_878), .C (n_776), .D (n_644), .Q
       (n_835));
  INX1 g92309(.A (n_732), .Q (n_834));
  NO2X1 g50573(.A (n_780), .B (n_708), .Q (n_833));
  NA3X1 g49821(.A (n_643), .B (n_642), .C (n_641), .Q (n_832));
  INX1 g92310(.A (n_8677), .Q (n_831));
  AND2X1 g92311(.A (n_944), .B (n_8162), .Q (n_830));
  ON22X1 g50396(.A (n_640), .B (alu_2nd_operand[2]), .C (n_693), .D
       (n_8496), .Q (n_829));
  NA2X1 g92312(.A (n_683), .B (n_6121), .Q (n_827));
  INX1 g92313(.A (n_6123), .Q (n_826));
  OA211X1 g50639(.A (n_687), .B (n_639), .C (n_638), .D (n_637), .Q
       (n_825));
  MU2IX1 g92314(.S (n_683), .IN0 (n_6134), .IN1 (\rs1_data[30]_39526 ),
       .Q (n_824));
  NA2X1 g92315(.A (alu_2nd_operand[2]), .B (n_828), .Q (n_823));
  ON221X1 g49729(.A (n_813), .B (n_897), .C (n_878), .D (n_895), .E
       (n_636), .Q (n_822));
  NO2X1 g49947(.A (n_635), .B (n_831), .Q (n_821));
  NA2X1 g49853(.A (n_634), .B (n_151), .Q (n_820));
  NO2X1 g92316(.A (n_831), .B (alu_2nd_operand[3]), .Q (n_819));
  MU2X1 g50397(.S (alu_2nd_operand[2]), .IN0 (n_633), .IN1 (n_632), .Q
       (n_818));
  OA222X1 g50577(.A (n_828), .B (n_698), .C (n_631), .D (n_166), .E
       (n_630), .F (n_826), .Q (n_817));
  NO2X1 g92317(.A (alu_2nd_operand[3]), .B (n_8677), .Q (n_816));
  AND4X1 g50638(.A (n_629), .B (n_628), .C (n_627), .D (n_626), .Q
       (n_815));
  AND4X1 g50643(.A (n_625), .B (n_624), .C (n_623), .D (n_622), .Q
       (n_814));
  INX1 g50503(.A (n_839), .Q (n_813));
  AND4X1 g50660(.A (n_621), .B (n_620), .C (n_619), .D (n_618), .Q
       (n_812));
  AN221X1 g49792(.A (read_data[27]), .B (n_617), .C (read_data[11]), .D
       (n_805), .E (n_616), .Q (n_811));
  ON22X1 g50313(.A (n_615), .B (n_898), .C (n_614), .D (n_896), .Q
       (n_810));
  ON211X1 g49722(.A (n_645), .B (n_776), .C (n_613), .D (n_612), .Q
       (n_809));
  MU2IX1 g50317(.S (alu_2nd_operand[2]), .IN0 (n_783), .IN1 (n_782), .Q
       (n_808));
  ON222X1 g49949(.A (n_898), .B (n_611), .C (n_173), .D (n_610), .E
       (n_609), .F (n_896), .Q (n_807));
  ON222X1 g49905(.A (n_153), .B (n_784), .C (n_776), .D (n_775), .E
       (n_781), .F (n_608), .Q (n_806));
  NO2X1 g92318(.A (n_607), .B (n_8073), .Q (n_805));
  AO221X1 g49824(.A (read_data[29]), .B (n_617), .C
       (\rs1_data[13]_39536 ), .D (n_606), .E (n_605), .Q (n_804));
  AO21X1 g49830(.A (n_604), .B (n_819), .C (n_820), .Q (n_803));
  ON222X1 g49950(.A (n_898), .B (n_603), .C (n_173), .D (n_602), .E
       (n_640), .F (n_896), .Q (n_802));
  MU2IX1 g50318(.S (alu_2nd_operand[2]), .IN0 (n_895), .IN1 (n_825), .Q
       (n_801));
  ON321X1 g49907(.A (n_708), .B (n_824), .C (n_601), .D (n_153), .E
       (n_897), .F (n_600), .Q (n_800));
  AO221X1 g49773(.A (read_data[14]), .B (n_805), .C (n_617), .D
       (read_data[30]), .E (n_599), .Q (n_799));
  MU2IX1 g50321(.S (alu_2nd_operand[2]), .IN0 (n_598), .IN1 (n_633), .Q
       (n_798));
  MU2IX1 g50238(.S (alu_2nd_operand[2]), .IN0 (n_632), .IN1 (n_817), .Q
       (n_797));
  MU2IX1 g50322(.S (alu_2nd_operand[2]), .IN0 (n_814), .IN1 (n_812), .Q
       (n_796));
  ON221X1 g49686(.A (n_813), .B (n_867), .C (n_878), .D (n_866), .E
       (n_597), .Q (n_795));
  NA2X1 g50591(.A (n_831), .B (n_914), .Q (n_794));
  MU2X1 g50390(.S (alu_2nd_operand[2]), .IN0 (n_614), .IN1 (n_169), .Q
       (n_793));
  NA2X1 g50574(.A (n_740), .B (n_830), .Q (n_792));
  AN21X1 g49764(.A (n_596), .B (n_595), .C (n_594), .Q (n_791));
  INX1 g49878(.A (n_593), .Q (n_790));
  NA2X1 g92319(.A (n_7264), .B (n_8296), .Q (n_789));
  OA211X1 g49760(.A (n_592), .B (n_170), .C (n_591), .D (n_590), .Q
       (n_788));
  NA2X1 g92320(.A (n_7263), .B (n_8296), .Q (n_787));
  OA211X1 g49743(.A (n_980), .B (n_794), .C (n_587), .D (n_586), .Q
       (n_786));
  NA2X1 g92321(.A (n_7262), .B (n_8296), .Q (n_785));
  AND4X1 g50646(.A (n_585), .B (n_584), .C (n_583), .D (n_582), .Q
       (n_784));
  AND4X1 g50645(.A (n_581), .B (n_580), .C (n_579), .D (n_578), .Q
       (n_783));
  AN211X1 g50640(.A (n_577), .B (n_6161), .C (n_576), .D (n_575), .Q
       (n_782));
  OA222X1 g92322(.A (n_639), .B (n_166), .C (n_828), .D (n_864), .E
       (n_630), .F (n_686), .Q (n_781));
  NA2X1 g92323(.A (n_574), .B (alu_2nd_operand[1]), .Q (n_780));
  MU2IX1 g92324(.S (alu_2nd_operand[0]), .IN0 (n_6181), .IN1 (n_6178),
       .Q (n_779));
  NA2X1 g92325(.A (n_577), .B (n_574), .Q (n_778));
  NA2X1 g92326(.A (n_828), .B (n_6167), .Q (n_777));
  NA2X2 g50593(.A (n_574), .B (n_914), .Q (n_776));
  AND4X1 g50665(.A (n_573), .B (n_572), .C (n_571), .D (n_570), .Q
       (n_775));
  OA22X1 g50181(.A (n_700), .B (n_813), .C (n_569), .D (n_153), .Q
       (n_774));
  INX1 g92327(.A (n_568), .Q (n_773));
  AN321X1 g49768(.A (n_830), .B (n_567), .C (n_165), .D (read_data[9]),
       .E (n_566), .F (n_565), .Q (n_772));
  AN221X1 g49767(.A (read_data[25]), .B (n_564), .C (read_data[17]), .D
       (n_697), .E (n_563), .Q (n_771));
  ON211X1 g49693(.A (n_977), .B (n_794), .C (n_562), .D (n_586), .Q
       (n_770));
  NA2X1 g92328(.A (n_7260), .B (n_8296), .Q (n_769));
  AN221X1 g49752(.A (n_830), .B (n_561), .C (n_922), .D (n_875), .E
       (n_560), .Q (n_768));
  NA3X1 g49692(.A (n_559), .B (n_558), .C (n_557), .Q (n_767));
  NA3X1 g49762(.A (n_556), .B (n_555), .C (n_554), .Q (n_766));
  NA2X1 g92329(.A (n_7257), .B (n_8296), .Q (n_765));
  OA211X1 g49802(.A (n_859), .B (n_725), .C (n_553), .D (n_552), .Q
       (n_764));
  AN211X1 g49779(.A (n_840), .B (n_936), .C (n_551), .D (n_550), .Q
       (n_763));
  NA2X1 g92330(.A (n_7256), .B (n_8296), .Q (n_762));
  AN21X1 g49801(.A (n_856), .B (n_549), .C (n_548), .Q (n_761));
  AN211X1 g49776(.A (n_915), .B (n_936), .C (n_547), .D (n_546), .Q
       (n_760));
  AN21X1 g49798(.A (n_1014), .B (n_549), .C (n_545), .Q (n_759));
  NA2X1 g92331(.A (n_7255), .B (n_8296), .Q (n_758));
  AND5X1 g49780(.A (n_544), .B (n_543), .C (n_542), .D (n_541), .E
       (n_540), .Q (n_757));
  NA2X1 g92332(.A (n_7254), .B (n_8296), .Q (n_756));
  AN21X1 g49800(.A (n_937), .B (n_549), .C (n_550), .Q (n_755));
  AN211X1 g49777(.A (n_938), .B (n_936), .C (n_539), .D (n_538), .Q
       (n_754));
  NO2X1 g49742(.A (n_537), .B (n_536), .Q (n_753));
  NA2X1 g92333(.A (n_7253), .B (n_8296), .Q (n_752));
  AN221X1 g49807(.A (n_740), .B (n_535), .C (n_8677), .D (n_807), .E
       (n_534), .Q (n_751));
  NA2X1 g92334(.A (n_7252), .B (n_8296), .Q (n_750));
  NA2X1 g92335(.A (n_531), .B (n_6149), .Q (n_748));
  NA2X1 g92336(.A (n_530), .B (\rs1_data[21]_39616 ), .Q (n_747));
  NA2X1 g92337(.A (n_164), .B (n_6141), .Q (n_746));
  NA2X1 g92338(.A (n_577), .B (\rs1_data[19]_39596 ), .Q (n_745));
  NA2X1 g92339(.A (n_531), .B (n_6145), .Q (n_744));
  NA2X1 g92340(.A (n_164), .B (n_6159), .Q (n_743));
  NA2X1 g92341(.A (n_530), .B (\rs1_data[25]_39346 ), .Q (n_742));
  NA2X1 g92342(.A (n_577), .B (n_6143), .Q (n_741));
  AND2X2 g92343(.A (n_831), .B (alu_2nd_operand[3]), .Q (n_740));
  NA3X1 g50629(.A (n_529), .B (n_528), .C (n_527), .Q (n_739));
  NA3X1 g50658(.A (n_526), .B (n_525), .C (n_524), .Q (n_738));
  AN221X1 g49774(.A (read_data[26]), .B (n_564), .C (read_data[18]), .D
       (n_697), .E (n_565), .Q (n_737));
  NA2X1 g92344(.A (n_566), .B (read_data[10]), .Q (n_736));
  AN211X1 g49822(.A (n_7280), .B (n_8296), .C (n_523), .D (n_522), .Q
       (n_735));
  NA2X1 g50592(.A (n_574), .B (n_830), .Q (n_734));
  NA2X1 g50576(.A (n_165), .B (n_914), .Q (n_733));
  MU2IX1 g92345(.S (alu_2nd_operand[0]), .IN0 (n_6123), .IN1 (n_6181),
       .Q (n_732));
  AND4X1 g50642(.A (n_521), .B (n_520), .C (n_519), .D (n_518), .Q
       (n_731));
  INX1 g50494(.A (n_833), .Q (n_730));
  MU2IX1 g92346(.S (alu_2nd_operand[0]), .IN0 (n_6178), .IN1 (n_6170),
       .Q (n_729));
  OA211X1 g49741(.A (n_517), .B (n_170), .C (n_533), .D (n_163), .Q
       (n_728));
  NA2X1 g92347(.A (n_7250), .B (n_8296), .Q (n_727));
  OA221X1 g49842(.A (n_648), .B (n_516), .C (n_515), .D (n_514), .E
       (n_513), .Q (n_726));
  NA2X1 g50583(.A (n_8677), .B (n_830), .Q (n_725));
  AN21X1 g49734(.A (n_7251), .B (n_8296), .C (n_512), .Q (n_724));
  AN21X1 g49786(.A (n_7279), .B (n_8296), .C (n_511), .Q (n_723));
  AN21X1 g50338(.A (n_911), .B (read_data[3]), .C (n_510), .Q (n_722));
  MU2IX1 g92348(.S (alu_2nd_operand[0]), .IN0 (n_6170), .IN1 (n_6165),
       .Q (n_721));
  AND4X1 g50644(.A (n_509), .B (n_508), .C (n_507), .D (n_506), .Q
       (n_720));
  AND4X1 g50633(.A (n_505), .B (n_504), .C (n_503), .D (n_502), .Q
       (n_719));
  OA211X1 g50641(.A (n_630), .B (n_501), .C (n_500), .D (n_499), .Q
       (n_718));
  OA222X1 g50578(.A (n_828), .B (n_824), .C (n_498), .D (n_166), .E
       (n_630), .F (n_639), .Q (n_717));
  NA2X1 g50519(.A (n_911), .B (read_data[4]), .Q (n_716));
  AN21X1 g49769(.A (n_7278), .B (n_8296), .C (n_495), .Q (n_715));
  AN222X1 g50523(.A (n_564), .B (read_data[28]), .C (read_data[12]), .D
       (n_566), .E (read_data[20]), .F (n_697), .Q (n_714));
  NA2X1 g92349(.A (n_531), .B (n_6139), .Q (n_713));
  NA2X1 g92350(.A (n_162), .B (n_6127), .Q (n_712));
  NA2X1 g92351(.A (n_530), .B (\rs1_data[11]_39506 ), .Q (n_711));
  NA2X1 g92352(.A (n_577), .B (n_6137), .Q (n_710));
  NA2X1 g92353(.A (n_740), .B (alu_2nd_operand[2]), .Q (n_709));
  INX1 g50671(.A (n_914), .Q (n_708));
  NA2X1 g92354(.A (n_531), .B (n_6141), .Q (n_707));
  NA2X1 g92355(.A (n_530), .B (\rs1_data[19]_39596 ), .Q (n_706));
  NA2X1 g92356(.A (n_164), .B (n_6132), .Q (n_705));
  NA2X1 g92357(.A (n_577), .B (n_8366), .Q (n_704));
  INX1 g50505(.A (n_776), .Q (n_703));
  NO2X1 g50331(.A (n_645), .B (n_813), .Q (n_702));
  INX1 g50245(.A (n_808), .Q (n_701));
  AND4X1 g50657(.A (n_493), .B (n_492), .C (n_491), .D (n_490), .Q
       (n_700));
  OA22X1 g50178(.A (n_775), .B (n_813), .C (n_569), .D (n_776), .Q
       (n_699));
  INX1 g92358(.A (n_567), .Q (n_698));
  ON21X1 g92359(.A (n_7708), .B (n_568), .C (n_487), .Q (n_697));
  AO221X1 g49756(.A (read_data[13]), .B (n_566), .C (n_564), .D
       (read_data[29]), .E (n_486), .Q (n_696));
  INX1 g50246(.A (n_801), .Q (n_695));
  AN22X1 g50183(.A (n_738), .B (n_839), .C (n_739), .D (n_837), .Q
       (n_694));
  AN221X1 g92360(.A (n_6178), .B (n_531), .C (n_6181), .D (n_530), .E
       (n_485), .Q (n_693));
  AO221X1 g49755(.A (read_data[14]), .B (n_566), .C (n_564), .D
       (read_data[30]), .E (n_484), .Q (n_692));
  NA2X1 g92361(.A (n_531), .B (\rs1_data[25]_39346 ), .Q (n_691));
  NA2X1 g92362(.A (n_577), .B (n_6145), .Q (n_690));
  NA2X1 g92363(.A (n_530), .B (n_6161), .Q (n_689));
  NA2X1 g92364(.A (n_162), .B (n_6143), .Q (n_688));
  INX1 g92365(.A (n_530), .Q (n_687));
  INX1 g92366(.A (\rs1_data[30]_39526 ), .Q (n_686));
  AN22X1 g92367(.A (n_164), .B (n_6135), .C (n_577), .D (n_6136), .Q
       (n_685));
  NA2X1 g92368(.A (n_531), .B (\rs1_data[29]_39416 ), .Q (n_684));
  INX2 g51948(.A (alu_2nd_operand[0]), .Q (n_683));
  ON22X1 g50177(.A (n_720), .B (n_776), .C (n_815), .D (n_153), .Q
       (n_682));
  AO221X1 g49757(.A (read_data[7]), .B (n_805), .C (n_617), .D
       (read_data[23]), .E (n_481), .Q (n_680));
  ON22X1 g50171(.A (n_879), .B (n_776), .C (n_645), .D (n_153), .Q
       (n_679));
  AO221X1 g49766(.A (read_data[8]), .B (n_805), .C (n_617), .D
       (read_data[24]), .E (n_480), .Q (n_678));
  INX1 g50323(.A (n_479), .Q (n_677));
  AN221X1 g49790(.A (read_data[25]), .B (n_617), .C (read_data[9]), .D
       (n_805), .E (n_478), .Q (n_676));
  NA2I1X1 g92371(.B (n_6134), .AN (alu_2nd_operand[31]), .Q (n_674));
  INX1 g92372(.A (n_477), .Q (n_673));
  ON22X1 g92373(.A (n_476), .B (n_843), .C (alu_2nd_operand[17]), .D
       (n_651), .Q (n_672));
  ON22X1 g92374(.A (alu_2nd_operand[19]), .B (n_475), .C
       (alu_2nd_operand[18]), .D (n_650), .Q (n_671));
  NA2X1 g92375(.A (alu_2nd_operand[19]), .B (n_475), .Q (n_670));
  NO2X1 g92376(.A (n_849), .B (n_474), .Q (n_669));
  NO2I1X1 g92377(.B (n_473), .AN (n_150), .Q (n_668));
  NO2X1 g92378(.A (n_472), .B (n_471), .Q (n_667));
  AN21X1 g92379(.A (n_8317), .B (n_686), .C (n_477), .Q (n_666));
  NO2X1 g92380(.A (n_470), .B (n_469), .Q (n_665));
  ON21X1 g92381(.A (n_468), .B (n_467), .C (n_466), .Q (n_664));
  NO2I1X1 g92382(.B (n_465), .AN (n_661), .Q (n_663));
  AO21X1 g92383(.A (n_464), .B (n_6135), .C (n_463), .Q (n_662));
  NA2X1 g92384(.A (alu_2nd_operand[27]), .B (n_462), .Q (n_661));
  ON21X1 g92385(.A (alu_2nd_operand[29]), .B (n_639), .C (n_461), .Q
       (n_660));
  ON21X1 g92386(.A (n_8317), .B (n_686), .C (n_674), .Q (n_659));
  ON21X1 g50537(.A (n_460), .B (n_459), .C (n_458), .Q (n_658));
  ON221X1 g49725(.A (n_457), .B (n_456), .C (n_455), .D (n_454), .E
       (n_453), .Q (n_657));
  AN21X1 g92387(.A (alu_2nd_operand[14]), .B (n_452), .C (n_451), .Q
       (n_656));
  AN21X1 g92388(.A (alu_2nd_operand[12]), .B (n_450), .C (n_449), .Q
       (n_655));
  ON32X1 g92389(.A (n_450), .B (alu_2nd_operand[12]), .C (n_449), .D
       (n_448), .E (alu_2nd_operand[13]), .Q (n_654));
  ON22X1 g92390(.A (alu_2nd_operand[15]), .B (n_447), .C
       (alu_2nd_operand[14]), .D (n_452), .Q (n_653));
  NA2X1 g92391(.A (alu_2nd_operand[15]), .B (n_447), .Q (n_652));
  INX1 g92392(.A (n_8366), .Q (n_651));
  INX1 g92393(.A (n_6141), .Q (n_650));
  INX1 g92394(.A (n_670), .Q (n_649));
  NA2X1 g92395(.A (n_740), .B (n_8496), .Q (n_648));
  NA2X1 g92396(.A (n_531), .B (n_6165), .Q (n_647));
  NA2X1 g92397(.A (n_530), .B (n_6183), .Q (n_646));
  AND4X1 g50666(.A (n_446), .B (n_445), .C (n_444), .D (n_443), .Q
       (n_645));
  OA21X1 g92398(.A (n_827), .B (alu_2nd_operand[1]), .C (n_152), .Q
       (n_644));
  AN22X1 g50194(.A (n_165), .B (n_442), .C (n_566), .D (read_data[8]),
       .Q (n_643));
  AN221X1 g49912(.A (n_1013), .B (n_7731), .C (read_data[16]), .D
       (n_697), .E (n_441), .Q (n_642));
  AN211X1 g49844(.A (n_564), .B (read_data[24]), .C (n_440), .D
       (n_439), .Q (n_641));
  AND4X1 g50653(.A (n_438), .B (n_519), .C (n_646), .D (n_710), .Q
       (n_640));
  NO2X4 g92399(.A (alu_2nd_operand[1]), .B (alu_2nd_operand[0]), .Q
       (n_164));
  INX1 g92400(.A (\rs1_data[29]_39416 ), .Q (n_639));
  AN22X1 g92401(.A (n_164), .B (n_6161), .C (n_577), .D (n_6135), .Q
       (n_638));
  NA2X1 g92402(.A (n_531), .B (n_6136), .Q (n_637));
  AN221X1 g49771(.A (read_data[26]), .B (n_617), .C (read_data[10]), .D
       (n_805), .E (n_437), .Q (n_636));
  OR2X1 g50244(.A (n_896), .B (n_436), .Q (n_635));
  NA3X1 g92403(.A (n_8623), .B (n_852), .C (n_8163), .Q (n_634));
  AND4X1 g50631(.A (n_628), .B (n_508), .C (n_435), .D (n_490), .Q
       (n_633));
  OA211X1 g50630(.A (n_630), .B (n_434), .C (n_433), .D (n_509), .Q
       (n_632));
  INX1 g92404(.A (n_6181), .Q (n_631));
  OR2X4 g92405(.A (alu_2nd_operand[1]), .B (n_683), .Q (n_630));
  NA2X1 g92406(.A (n_531), .B (\rs1_data[13]_39536 ), .Q (n_629));
  NA2X1 g92407(.A (n_164), .B (\rs1_data[11]_39506 ), .Q (n_628));
  NA2X1 g92408(.A (n_530), .B (n_6153), .Q (n_627));
  NA2X1 g92409(.A (n_577), .B (\rs1_data[12]_39516 ), .Q (n_626));
  NA2X1 g92410(.A (n_531), .B (n_8366), .Q (n_625));
  NA2X1 g92411(.A (n_530), .B (n_6141), .Q (n_624));
  NA2X1 g92412(.A (n_164), .B (n_6155), .Q (n_623));
  NA2X1 g92413(.A (n_577), .B (n_6132), .Q (n_622));
  NA2X1 g92414(.A (n_531), .B (\rs1_data[21]_39616 ), .Q (n_621));
  NA2X1 g92415(.A (n_164), .B (\rs1_data[19]_39596 ), .Q (n_620));
  NA2X1 g92416(.A (n_530), .B (n_6159), .Q (n_619));
  NA2X1 g92417(.A (n_577), .B (n_6149), .Q (n_618));
  AND3X1 g92418(.A (n_8566), .B (n_852), .C (n_7303), .Q (n_617));
  ON221X1 g49862(.A (n_432), .B (n_431), .C (n_430), .D (n_429), .E
       (n_428), .Q (n_616));
  AND4X1 g50664(.A (n_521), .B (n_713), .C (n_528), .D (n_446), .Q
       (n_615));
  AND4X1 g50651(.A (n_647), .B (n_712), .C (n_520), .D (n_427), .Q
       (n_614));
  OA22X1 g50182(.A (n_877), .B (n_153), .C (n_717), .D (n_608), .Q
       (n_613));
  AN221X1 g49772(.A (read_data[28]), .B (n_617), .C (read_data[12]), .D
       (n_805), .E (n_426), .Q (n_612));
  AND4X1 g50663(.A (n_491), .B (n_507), .C (n_626), .D (n_570), .Q
       (n_611));
  INX1 g50326(.A (n_873), .Q (n_610));
  AND4X1 g50655(.A (n_492), .B (n_425), .C (n_506), .D (n_424), .Q
       (n_609));
  OR2X1 g50566(.A (n_149), .B (n_708), .Q (n_608));
  AN21X1 g92419(.A (n_957), .B (n_7303), .C (n_8487), .Q (n_607));
  ON211X1 g50206(.A (alu_2nd_operand[13]), .B (n_432), .C (n_430), .D
       (n_423), .Q (n_606));
  ON221X1 g50200(.A (n_432), .B (n_422), .C (n_430), .D (n_421), .E
       (n_420), .Q (n_605));
  NO2X1 g50243(.A (n_167), .B (n_436), .Q (n_604));
  AND4X1 g50662(.A (n_419), .B (n_711), .C (n_443), .D (n_418), .Q
       (n_603));
  INX1 g50327(.A (n_869), .Q (n_602));
  NA2X1 g92420(.A (n_167), .B (n_819), .Q (n_601));
  NA2X1 g50335(.A (n_738), .B (n_703), .Q (n_600));
  AO221X1 g49827(.A (n_6153), .B (n_417), .C (alu_2nd_operand[14]), .D
       (n_416), .E (n_415), .Q (n_599));
  AND4X1 g50650(.A (n_629), .B (n_493), .C (n_623), .D (n_572), .Q
       (n_598));
  AN211X1 g49733(.A (n_805), .B (read_data[15]), .C (n_414), .D
       (n_413), .Q (n_597));
  INX1 g50596(.A (n_615), .Q (n_596));
  NO2X1 g50580(.A (n_494), .B (n_170), .Q (n_595));
  ON221X1 g49787(.A (n_734), .B (n_412), .C (n_411), .D (n_601), .E
       (n_410), .Q (n_594));
  NA2X2 g49962(.A (n_409), .B (n_408), .Q (n_593));
  AN21X1 g49886(.A (n_479), .B (n_740), .C (n_407), .Q (n_592));
  AN21X1 g49813(.A (n_406), .B (alu_2nd_operand[1]), .C (n_593), .Q
       (n_591));
  AN221X1 g49867(.A (n_405), .B (n_843), .C (n_404), .D (n_8366), .E
       (n_403), .Q (n_590));
  AN21X1 g49880(.A (n_829), .B (n_740), .C (n_402), .Q (n_589));
  AND3X1 g49782(.A (n_591), .B (n_401), .C (n_400), .Q (n_588));
  AN21X1 g49775(.A (n_399), .B (n_830), .C (n_398), .Q (n_587));
  NO2X1 g49849(.A (n_593), .B (n_406), .Q (n_586));
  NA2X1 g92421(.A (n_530), .B (n_6149), .Q (n_585));
  NA2X1 g92422(.A (n_531), .B (\rs1_data[19]_39596 ), .Q (n_584));
  NA2X1 g92423(.A (n_577), .B (n_6141), .Q (n_583));
  NA2X1 g92424(.A (n_164), .B (n_8366), .Q (n_582));
  NA2X1 g92425(.A (n_530), .B (n_6145), .Q (n_581));
  NA2X1 g92426(.A (n_577), .B (n_6159), .Q (n_580));
  NA2X1 g92427(.A (n_531), .B (n_6143), .Q (n_579));
  NA2X1 g92428(.A (n_164), .B (\rs1_data[21]_39616 ), .Q (n_578));
  INX4 g92429(.A (n_630), .Q (n_577));
  INX1 g92430(.A (n_397), .Q (n_576));
  ON21X1 g92431(.A (n_489), .B (n_462), .C (n_396), .Q (n_575));
  NO2X1 g92432(.A (n_898), .B (n_8677), .Q (n_574));
  NA2X1 g92433(.A (n_530), .B (n_6132), .Q (n_573));
  NA2X1 g92434(.A (n_577), .B (n_6153), .Q (n_572));
  NA2X1 g92435(.A (n_531), .B (n_6155), .Q (n_571));
  NA2X1 g92436(.A (n_164), .B (\rs1_data[13]_39536 ), .Q (n_570));
  OA211X1 g50565(.A (n_721), .B (alu_2nd_operand[1]), .C (n_435), .D
       (n_425), .Q (n_569));
  NA2X1 g92437(.A (n_852), .B (n_7302), .Q (n_568));
  ON21X1 g92438(.A (alu_2nd_operand[0]), .B (n_395), .C (n_394), .Q
       (n_567));
  NO2X1 g92439(.A (n_7710), .B (n_568), .Q (n_566));
  NO2X1 g49831(.A (n_393), .B (n_828), .Q (n_565));
  NO2X1 g92440(.A (n_7707), .B (n_568), .Q (n_564));
  AO211X1 g49826(.A (n_8566), .B (n_8296), .C (n_392), .D (n_391), .Q
       (n_563));
  AN221X1 g49748(.A (n_390), .B (n_881), .C (n_882), .D (n_389), .E
       (n_388), .Q (n_562));
  ON221X1 g49903(.A (n_648), .B (n_611), .C (n_709), .D (n_609), .E
       (n_387), .Q (n_561));
  ON211X1 g49781(.A (n_386), .B (n_862), .C (n_557), .D (n_385), .Q
       (n_560));
  NA2X1 g49835(.A (n_871), .B (n_922), .Q (n_559));
  AN221X1 g49747(.A (n_390), .B (n_869), .C (n_882), .D (n_384), .E
       (n_383), .Q (n_558));
  AN21X1 g49850(.A (n_604), .B (n_740), .C (n_593), .Q (n_557));
  AN21X1 g49808(.A (n_798), .B (n_382), .C (n_381), .Q (n_556));
  AN221X1 g49811(.A (n_6143), .B (n_380), .C (n_922), .D (n_967), .E
       (n_379), .Q (n_555));
  INX2 g49834(.A (n_550), .Q (n_554));
  OA22X1 g50166(.A (n_412), .B (n_378), .C (n_615), .D (n_377), .Q
       (n_553));
  OA22X1 g50174(.A (n_376), .B (n_734), .C (n_375), .D (n_374), .Q
       (n_552));
  ON221X1 g49858(.A (n_432), .B (n_373), .C (n_430), .D (n_372), .E
       (n_371), .Q (n_551));
  NA2X2 g49854(.A (n_790), .B (n_370), .Q (n_550));
  INX1 g50499(.A (n_725), .Q (n_549));
  ON221X1 g49897(.A (n_374), .B (n_369), .C (n_377), .D (n_611), .E
       (n_368), .Q (n_548));
  ON221X1 g49864(.A (n_432), .B (n_367), .C (n_430), .D (n_366), .E
       (n_365), .Q (n_547));
  ON21X1 g49814(.A (n_635), .B (n_828), .C (n_554), .Q (n_546));
  ON221X1 g49896(.A (n_378), .B (n_364), .C (n_377), .D (n_603), .E
       (n_363), .Q (n_545));
  INX1 g49797(.A (n_546), .Q (n_544));
  NA2I1X1 g50163(.B (n_936), .AN (n_943), .Q (n_543));
  ON21X1 g50553(.A (n_465), .B (n_463), .C (n_405), .Q (n_542));
  ON21X1 g50525(.A (alu_2nd_operand[26]), .B (n_6161), .C (n_362), .Q
       (n_541));
  AN321X0 g50218(.A (n_6161), .B (n_361), .C (alu_2nd_operand[26]), .D
       (n_8157), .E (csr_data_out[26]), .F (n_360), .Q (n_540));
  ON221X1 g49856(.A (n_462), .B (n_359), .C (n_432), .D (n_661), .E
       (n_358), .Q (n_539));
  ON221X1 g49810(.A (n_374), .B (n_516), .C (n_377), .D (n_598), .E
       (n_357), .Q (n_538));
  ON21X1 g49761(.A (n_933), .B (n_725), .C (n_356), .Q (n_537));
  ON21X1 g49805(.A (n_355), .B (n_170), .C (n_554), .Q (n_536));
  MU2IX1 g50394(.S (alu_2nd_operand[2]), .IN0 (n_369), .IN1 (n_354), .Q
       (n_535));
  ON321X1 g50169(.A (n_639), .B (alu_2nd_operand[0]), .C (n_353), .D
       (n_352), .E (n_780), .F (n_351), .Q (n_534));
  NO2X1 g49812(.A (n_550), .B (n_604), .Q (n_533));
  AND2X4 g92441(.A (alu_2nd_operand[1]), .B (n_683), .Q (n_531));
  AND2X4 g92442(.A (alu_2nd_operand[1]), .B (alu_2nd_operand[0]), .Q
       (n_530));
  AND2X1 g92443(.A (n_438), .B (n_419), .Q (n_529));
  NA2X1 g92444(.A (n_577), .B (\rs1_data[11]_39506 ), .Q (n_528));
  NA2X1 g92445(.A (n_530), .B (\rs1_data[13]_39536 ), .Q (n_527));
  AND2X1 g92446(.A (n_349), .B (n_418), .Q (n_526));
  NA2X1 g92447(.A (n_530), .B (n_8366), .Q (n_525));
  NA2X1 g92448(.A (n_531), .B (n_6132), .Q (n_524));
  AN21X1 g50551(.A (n_348), .B (n_347), .C (n_432), .Q (n_523));
  ON311X1 g49914(.A (n_161), .B (n_826), .C (n_8496), .D (n_346), .E
       (n_345), .Q (n_522));
  NA2X1 g92449(.A (n_530), .B (n_6137), .Q (n_521));
  NA2X1 g92450(.A (n_577), .B (n_6183), .Q (n_520));
  NA2X1 g92451(.A (n_531), .B (n_6127), .Q (n_519));
  NA2X1 g92452(.A (n_164), .B (n_6165), .Q (n_518));
  AN221X1 g49804(.A (n_740), .B (n_384), .C (n_8677), .D (n_802), .E
       (n_344), .Q (n_517));
  AND4X1 g50649(.A (n_585), .B (n_621), .C (n_580), .D (n_688), .Q
       (n_516));
  INX1 g92453(.A (n_574), .Q (n_515));
  OA211X1 g50678(.A (n_864), .B (alu_2nd_operand[1]), .C (n_396), .D
       (n_684), .Q (n_514));
  OA222X1 g49906(.A (n_494), .B (n_8591), .C (n_686), .D (n_778), .E
       (n_340), .F (n_709), .Q (n_513));
  ON211X0 g49765(.A (n_733), .B (n_864), .C (n_339), .D (n_409), .Q
       (n_512));
  ON211X1 g49823(.A (n_338), .B (n_631), .C (n_393), .D (n_337), .Q
       (n_511));
  AO222X1 g50522(.A (read_data[27]), .B (n_564), .C (read_data[19]), .D
       (n_697), .E (read_data[11]), .F (n_566), .Q (n_510));
  NA2X1 g92454(.A (n_162), .B (n_6183), .Q (n_509));
  NA2X1 g92455(.A (n_531), .B (n_6137), .Q (n_508));
  NA2X1 g92456(.A (n_530), .B (n_6139), .Q (n_507));
  NA2X1 g92457(.A (n_577), .B (n_6127), .Q (n_506));
  NA2X1 g92458(.A (n_530), .B (n_6143), .Q (n_505));
  NA2X1 g92459(.A (n_531), .B (n_6159), .Q (n_504));
  NA2X1 g92460(.A (n_162), .B (n_6149), .Q (n_503));
  NA2X1 g92461(.A (n_577), .B (\rs1_data[21]_39616 ), .Q (n_502));
  AN21X1 g92463(.A (n_531), .B (n_6161), .C (n_336), .Q (n_500));
  NA2X1 g92464(.A (n_162), .B (n_6145), .Q (n_499));
  INX1 g92465(.A (n_6136), .Q (n_498));
  INX1 g92466(.A (n_6178), .Q (n_497));
  AN22X1 g92467(.A (n_531), .B (n_6123), .C (n_530), .D (n_6167), .Q
       (n_496));
  ON211X1 g49794(.A (n_335), .B (n_432), .C (n_334), .D (n_393), .Q
       (n_495));
  NA2X1 g92468(.A (n_816), .B (alu_2nd_operand[2]), .Q (n_494));
  NA2X1 g92469(.A (n_530), .B (\rs1_data[12]_39516 ), .Q (n_493));
  NA2X1 g92470(.A (n_162), .B (n_6137), .Q (n_492));
  NA2X1 g92471(.A (n_531), .B (\rs1_data[11]_39506 ), .Q (n_491));
  NA2X1 g92472(.A (n_577), .B (n_6139), .Q (n_490));
  INX1 g92473(.A (n_531), .Q (n_489));
  AN22X1 g92474(.A (n_164), .B (n_6170), .C (n_577), .D (n_6178), .Q
       (n_488));
  INX1 g92475(.A (n_617), .Q (n_487));
  ON211X1 g49795(.A (n_333), .B (n_432), .C (n_332), .D (n_331), .Q
       (n_486));
  ON21X1 g92476(.A (n_630), .B (n_330), .C (n_518), .Q (n_485));
  NA3X1 g49793(.A (n_332), .B (n_329), .C (n_328), .Q (n_484));
  NA3X1 g49796(.A (n_151), .B (n_323), .C (n_322), .Q (n_481));
  ON21X1 g49817(.A (n_321), .B (n_432), .C (n_320), .Q (n_480));
  MU2IX1 g50392(.S (alu_2nd_operand[2]), .IN0 (n_609), .IN1 (n_168), .Q
       (n_479));
  ON211X1 g49837(.A (n_319), .B (n_432), .C (n_318), .D (n_317), .Q
       (n_478));
  AND2X1 g92478(.A (alu_2nd_operand[31]), .B (n_316), .Q (n_477));
  INX1 g92479(.A (n_315), .Q (n_476));
  INX1 g92480(.A (\rs1_data[19]_39596 ), .Q (n_475));
  NA3X1 g92481(.A (n_663), .B (n_148), .C (n_314), .Q (n_474));
  AND2X1 g92482(.A (alu_2nd_operand[22]), .B (n_313), .Q (n_473));
  NO2I1X1 g92483(.B (n_6149), .AN (alu_2nd_operand[20]), .Q (n_472));
  NO2X1 g92484(.A (n_312), .B (\rs1_data[21]_39616 ), .Q (n_471));
  AND2X1 g92485(.A (alu_2nd_operand[28]), .B (n_498), .Q (n_470));
  INX1 g92486(.A (n_311), .Q (n_469));
  NA2I1X1 g92487(.B (n_6145), .AN (alu_2nd_operand[24]), .Q (n_468));
  INX1 g92488(.A (n_314), .Q (n_467));
  OR2X1 g92489(.A (alu_2nd_operand[25]), .B (n_501), .Q (n_466));
  AND2X1 g92490(.A (alu_2nd_operand[26]), .B (n_310), .Q (n_465));
  INX1 g92491(.A (alu_2nd_operand[27]), .Q (n_464));
  NO2X1 g92492(.A (alu_2nd_operand[26]), .B (n_310), .Q (n_463));
  INX1 g92493(.A (n_6135), .Q (n_462));
  NA2X1 g92494(.A (n_309), .B (n_311), .Q (n_461));
  AN22X1 g50886(.A (n_308), .B (n_307), .C (n_312), .D
       (\rs1_data[21]_39616 ), .Q (n_460));
  INX1 g92495(.A (n_668), .Q (n_459));
  ON21X1 g92496(.A (n_306), .B (n_305), .C (n_150), .Q (n_458));
  INX1 g92497(.A (n_304), .Q (n_457));
  OA21X1 g92498(.A (n_303), .B (n_321), .C (n_302), .Q (n_456));
  NO2I1X1 g92499(.B (\rs1_data[11]_39506 ), .AN (alu_2nd_operand[11]),
       .Q (n_455));
  AND2X1 g92500(.A (n_301), .B (n_300), .Q (n_454));
  ON311X1 g49749(.A (n_299), .B (n_298), .C (n_297), .D (n_304), .E
       (n_296), .Q (n_453));
  INX1 g51932(.A (n_6153), .Q (n_452));
  INX1 g92501(.A (n_652), .Q (n_451));
  INX1 g51933(.A (\rs1_data[12]_39516 ), .Q (n_450));
  INX1 g92502(.A (n_422), .Q (n_449));
  INX1 g92503(.A (\rs1_data[13]_39536 ), .Q (n_448));
  INX1 g92504(.A (n_6155), .Q (n_447));
  NA2X1 g92505(.A (n_164), .B (\rs1_data[12]_39516 ), .Q (n_446));
  NA2X1 g92506(.A (n_531), .B (n_6153), .Q (n_445));
  NA2X1 g92507(.A (n_530), .B (n_6155), .Q (n_444));
  NA2X1 g92508(.A (n_577), .B (\rs1_data[13]_39536 ), .Q (n_443));
  NO2X1 g50570(.A (n_827), .B (n_170), .Q (n_442));
  NO2X1 g50348(.A (n_853), .B (n_295), .Q (n_441));
  AN21X1 g50531(.A (n_827), .B (n_294), .C (n_432), .Q (n_440));
  ON221X1 g50202(.A (n_161), .B (n_394), .C (n_430), .D (n_293), .E
       (n_292), .Q (n_439));
  NA2X1 g92509(.A (n_162), .B (n_6139), .Q (n_438));
  ON21X1 g49819(.A (n_301), .B (n_432), .C (n_291), .Q (n_437));
  NA3X1 g50404(.A (n_6134), .B (n_914), .C (alu_operation_code_39112),
       .Q (n_436));
  NA2X1 g92510(.A (n_530), .B (n_6127), .Q (n_435));
  INX1 g51943(.A (n_6165), .Q (n_434));
  AN22X1 g92511(.A (n_531), .B (n_6170), .C (n_530), .D (n_6178), .Q
       (n_433));
  INX3 g50675(.A (n_405), .Q (n_432));
  NO2X1 g92512(.A (n_455), .B (n_290), .Q (n_431));
  INX3 g50674(.A (n_362), .Q (n_430));
  NO2X1 g92513(.A (alu_2nd_operand[11]), .B (\rs1_data[11]_39506 ), .Q
       (n_429));
  AN31X1 g50220(.A (n_361), .B (\rs1_data[11]_39506 ), .C
       (alu_2nd_operand[11]), .D (n_289), .Q (n_428));
  NA2X1 g92514(.A (n_530), .B (n_6170), .Q (n_427));
  AO221X1 g49818(.A (\rs1_data[12]_39516 ), .B (n_288), .C
       (alu_2nd_operand[12]), .D (n_287), .E (n_286), .Q (n_426));
  NA2X1 g92515(.A (n_531), .B (n_6183), .Q (n_425));
  NA2X1 g92516(.A (n_530), .B (n_6165), .Q (n_424));
  NA2X1 g50544(.A (alu_2nd_operand[13]), .B (n_361), .Q (n_423));
  NA2X1 g92517(.A (alu_2nd_operand[13]), .B (n_448), .Q (n_422));
  INX1 g92518(.A (alu_2nd_operand[13]), .Q (n_421));
  AN222X1 g92519(.A (n_8166), .B (n_7689), .C (n_7937), .D (n_2548), .E
       (csr_data_out[13]), .F (n_8157), .Q (n_420));
  NA2X1 g92520(.A (n_531), .B (\rs1_data[12]_39516 ), .Q (n_419));
  NA2X1 g92521(.A (n_162), .B (n_6153), .Q (n_418));
  ON21X1 g50356(.A (alu_2nd_operand[14]), .B (n_432), .C (n_430), .Q
       (n_417));
  ON221X1 g50226(.A (n_161), .B (n_452), .C (n_432), .D (n_6153), .E
       (n_430), .Q (n_416));
  AO222X1 g92522(.A (n_8166), .B (n_7688), .C (n_8157), .D
       (csr_data_out[14]), .E (n_7938), .F (n_2548), .Q (n_415));
  ON311X1 g49770(.A (n_708), .B (n_864), .C (n_601), .D (n_285), .E
       (n_284), .Q (n_414));
  INX1 g50670(.A (n_634), .Q (n_413));
  AND4X1 g50661(.A (n_705), .B (n_445), .C (n_527), .D (n_349), .Q
       (n_412));
  INX1 g50493(.A (n_442), .Q (n_411));
  AND3X1 g49863(.A (n_283), .B (n_282), .C (n_281), .Q (n_410));
  NO2X1 g50569(.A (n_413), .B (n_280), .Q (n_409));
  NA2X1 g50239(.A (n_8677), .B (n_279), .Q (n_408));
  ON222X1 g50167(.A (n_515), .B (n_354), .C (n_494), .D (n_611), .E
       (n_601), .F (n_698), .Q (n_407));
  NO2X1 g49953(.A (n_370), .B (n_8496), .Q (n_406));
  AND2X2 g92523(.A (n_944), .B (n_8161), .Q (n_405));
  ON211X1 g50224(.A (alu_2nd_operand[17]), .B (n_432), .C (n_430), .D
       (n_278), .Q (n_404));
  AO221X1 g50364(.A (n_362), .B (alu_2nd_operand[17]), .C (n_8157), .D
       (csr_data_out[17]), .E (n_277), .Q (n_403));
  ON222X1 g50168(.A (n_494), .B (n_603), .C (n_515), .D (n_364), .E
       (n_946), .F (n_149), .Q (n_402));
  NA2X1 g50222(.A (n_276), .B (n_6141), .Q (n_401));
  AN221X1 g49855(.A (n_8157), .B (csr_data_out[18]), .C
       (alu_2nd_operand[18]), .D (n_275), .E (n_274), .Q (n_400));
  ON222X1 g49904(.A (n_494), .B (n_598), .C (n_515), .D (n_340), .E
       (n_817), .F (n_149), .Q (n_399));
  ON21X1 g49809(.A (n_818), .B (n_792), .C (n_273), .Q (n_398));
  NA2X1 g92524(.A (n_162), .B (\rs1_data[25]_39346 ), .Q (n_397));
  NA2X1 g92525(.A (n_530), .B (n_6136), .Q (n_396));
  INX1 g92526(.A (n_6167), .Q (n_395));
  NA2X1 g92527(.A (alu_2nd_operand[0]), .B (n_6121), .Q (n_394));
  OR2X1 g49875(.A (n_151), .B (n_8496), .Q (n_393));
  AN21X1 g50558(.A (n_777), .B (n_272), .C (n_432), .Q (n_392));
  ON311X1 g49915(.A (n_161), .B (n_395), .C (n_828), .D (n_271), .E
       (n_270), .Q (n_391));
  INX1 g50496(.A (n_269), .Q (n_390));
  MU2IX1 g50391(.S (alu_2nd_operand[2]), .IN0 (n_375), .IN1 (n_412), .Q
       (n_389));
  ON221X1 g49783(.A (n_378), .B (n_615), .C (n_377), .D (n_614), .E
       (n_268), .Q (n_388));
  NA2X1 g50179(.A (n_873), .B (n_819), .Q (n_387));
  INX1 g50324(.A (n_535), .Q (n_386));
  AN221X1 g49861(.A (n_405), .B (n_471), .C (n_267), .D
       (\rs1_data[21]_39616 ), .E (n_266), .Q (n_385));
  MU2IX1 g50315(.S (alu_2nd_operand[2]), .IN0 (n_265), .IN1 (n_364), .Q
       (n_384));
  ON221X1 g49784(.A (n_378), .B (n_603), .C (n_377), .D (n_640), .E
       (n_264), .Q (n_383));
  INX1 g50495(.A (n_792), .Q (n_382));
  ON222X1 g49841(.A (n_734), .B (n_516), .C (n_269), .D (n_863), .E
       (n_340), .F (n_374), .Q (n_381));
  ON211X1 g50210(.A (alu_2nd_operand[23]), .B (n_432), .C (n_430), .D
       (n_263), .Q (n_380));
  ON21X1 g50203(.A (n_150), .B (n_432), .C (n_262), .Q (n_379));
  OR2X1 g50582(.A (n_648), .B (n_170), .Q (n_378));
  OR2X1 g50581(.A (n_709), .B (n_170), .Q (n_377));
  AND4X1 g50632(.A (n_504), .B (n_747), .C (n_499), .D (n_741), .Q
       (n_376));
  AND4X1 g50635(.A (n_707), .B (n_525), .C (n_503), .D (n_745), .Q
       (n_375));
  INX1 g50498(.A (n_595), .Q (n_374));
  AND2X1 g92528(.A (n_468), .B (n_148), .Q (n_373));
  NO2X1 g92529(.A (alu_2nd_operand[24]), .B (n_6145), .Q (n_372));
  AN321X1 g50217(.A (n_6145), .B (n_361), .C (alu_2nd_operand[24]), .D
       (n_8157), .E (csr_data_out[24]), .F (n_261), .Q (n_371));
  NA2X1 g50236(.A (alu_2nd_operand[3]), .B (n_279), .Q (n_370));
  AND4X1 g50636(.A (n_584), .B (n_624), .C (n_578), .D (n_618), .Q
       (n_369));
  OA22X1 g50173(.A (n_260), .B (n_734), .C (n_354), .D (n_378), .Q
       (n_368));
  AND2X1 g92530(.A (n_466), .B (n_314), .Q (n_367));
  NO2X1 g92531(.A (alu_2nd_operand[25]), .B (\rs1_data[25]_39346 ), .Q
       (n_366));
  AN321X1 g50223(.A (\rs1_data[25]_39346 ), .B (n_361), .C
       (alu_2nd_operand[25]), .D (n_8157), .E (csr_data_out[25]), .F
       (n_259), .Q (n_365));
  AND4X1 g50654(.A (n_746), .B (n_524), .C (n_444), .D (n_704), .Q
       (n_364));
  OA22X1 g50175(.A (n_265), .B (n_374), .C (n_258), .D (n_734), .Q
       (n_363));
  AND2X2 g92532(.A (n_944), .B (n_8159), .Q (n_362));
  AND2X2 g92533(.A (n_944), .B (n_8158), .Q (n_361));
  AO222X1 g92534(.A (read_data[26]), .B (n_160), .C (n_8166), .D
       (n_7675), .E (n_7951), .F (n_2548), .Q (n_360));
  AN211X1 g50205(.A (alu_2nd_operand[27]), .B (n_361), .C (n_362), .D
       (n_257), .Q (n_359));
  AN221X1 g50358(.A (n_8157), .B (csr_data_out[27]), .C
       (alu_2nd_operand[27]), .D (n_362), .E (n_256), .Q (n_358));
  OA211X1 g49788(.A (n_717), .B (n_776), .C (n_635), .D (n_255), .Q
       (n_356));
  AN21X1 g49889(.A (n_389), .B (n_740), .C (n_254), .Q (n_355));
  AND4X1 g50659(.A (n_582), .B (n_571), .C (n_627), .D (n_622), .Q
       (n_354));
  INX1 g92535(.A (n_165), .Q (n_353));
  MU2IX1 g92536(.S (alu_2nd_operand[0]), .IN0 (n_6135), .IN1 (n_6161),
       .Q (n_352));
  OA22X1 g50332(.A (n_260), .B (n_494), .C (n_778), .D (n_498), .Q
       (n_351));
  AN221X1 g49860(.A (n_405), .B (n_469), .C (n_253), .D
       (\rs1_data[29]_39416 ), .E (n_252), .Q (n_350));
  NA2X1 g92537(.A (n_577), .B (n_6155), .Q (n_349));
  NA2X1 g92538(.A (n_8496), .B (n_6123), .Q (n_348));
  NA2X1 g92539(.A (alu_2nd_operand[2]), .B (n_826), .Q (n_347));
  AN222X1 g92540(.A (n_8157), .B (csr_data_out[2]), .C (n_7925), .D
       (n_2548), .E (n_7681), .F (n_8166), .Q (n_346));
  ON21X1 g50564(.A (alu_2nd_operand[2]), .B (n_6123), .C (n_362), .Q
       (n_345));
  ON222X1 g49909(.A (n_515), .B (n_251), .C (n_494), .D (n_258), .E
       (n_778), .F (n_639), .Q (n_344));
  OA21X1 g50355(.A (n_8317), .B (n_432), .C (n_430), .Q (n_343));
  AN221X1 g49869(.A (n_8157), .B (csr_data_out[30]), .C (n_8317), .D
       (n_250), .E (n_249), .Q (n_342));
  AND4X1 g50669(.A (n_573), .B (n_620), .C (n_625), .D (n_583), .Q
       (n_340));
  OA211X1 g49825(.A (n_853), .B (n_432), .C (n_246), .D (n_245), .Q
       (n_339));
  AN221X1 g50204(.A (n_405), .B (n_173), .C (n_361), .D
       (alu_2nd_operand[3]), .E (n_362), .Q (n_338));
  AN221X1 g50201(.A (n_362), .B (alu_2nd_operand[3]), .C (n_405), .D
       (n_244), .E (n_243), .Q (n_337));
  INX1 g92541(.A (n_242), .Q (n_336));
  NA2X1 g92542(.A (n_831), .B (n_6178), .Q (n_335));
  AN221X1 g49872(.A (n_362), .B (n_6178), .C (n_241), .D (n_8677), .E
       (n_240), .Q (n_334));
  OR2X1 g92543(.A (alu_2nd_operand[5]), .B (n_330), .Q (n_333));
  OR2X1 g49874(.A (n_151), .B (n_167), .Q (n_332));
  AN221X1 g49866(.A (n_362), .B (n_6170), .C (n_239), .D
       (alu_2nd_operand[5]), .E (n_238), .Q (n_331));
  INX1 g92544(.A (n_6170), .Q (n_330));
  NA2X1 g50557(.A (n_298), .B (n_405), .Q (n_329));
  AN221X1 g49868(.A (n_362), .B (n_6165), .C (n_237), .D
       (alu_2nd_operand[6]), .E (n_236), .Q (n_328));
  AND2X1 g92545(.A (n_8165), .B (read_data[7]), .Q (n_327));
  NO2I1X2 g92546(.B (n_7710), .AN (read_data[15]), .Q (n_326));
  NO2I1X1 g92547(.B (n_7708), .AN (read_data[23]), .Q (n_325));
  NO2I1X1 g92548(.B (n_7707), .AN (read_data[31]), .Q (n_324));
  NA2X1 g50529(.A (n_299), .B (n_405), .Q (n_323));
  AN221X1 g49871(.A (n_362), .B (n_6183), .C (n_235), .D
       (alu_2nd_operand[7]), .E (n_234), .Q (n_322));
  OR2X1 g92549(.A (alu_2nd_operand[8]), .B (n_233), .Q (n_321));
  AN221X1 g49873(.A (n_362), .B (n_6127), .C (n_232), .D
       (alu_2nd_operand[8]), .E (n_231), .Q (n_320));
  NO2I1X1 g92550(.B (n_303), .AN (n_302), .Q (n_319));
  AN31X1 g50209(.A (n_361), .B (n_6137), .C (alu_2nd_operand[9]), .D
       (n_230), .Q (n_318));
  ON21X1 g50534(.A (alu_2nd_operand[9]), .B (n_6137), .C (n_362), .Q
       (n_317));
  INX1 g92551(.A (n_6134), .Q (n_316));
  NO2X1 g92552(.A (n_8495), .B (n_229), .Q (n_315));
  NA2X1 g92553(.A (alu_2nd_operand[25]), .B (n_501), .Q (n_314));
  INX1 g92554(.A (n_6159), .Q (n_313));
  INX1 g92555(.A (alu_2nd_operand[21]), .Q (n_312));
  NA2X1 g92556(.A (alu_2nd_operand[29]), .B (n_639), .Q (n_311));
  INX1 g92557(.A (n_6161), .Q (n_310));
  NO2X1 g92558(.A (alu_2nd_operand[28]), .B (n_498), .Q (n_309));
  NO2I1X1 g92559(.B (alu_2nd_operand[20]), .AN (n_6149), .Q (n_308));
  INX1 g92560(.A (n_471), .Q (n_307));
  NO2I1X1 g92561(.B (alu_2nd_operand[22]), .AN (n_6159), .Q (n_306));
  NO2I1X1 g92562(.B (alu_2nd_operand[23]), .AN (n_6143), .Q (n_305));
  AN21X1 g92563(.A (alu_2nd_operand[10]), .B (n_228), .C (n_455), .Q
       (n_304));
  NO2I1X1 g92564(.B (n_6137), .AN (alu_2nd_operand[9]), .Q (n_303));
  NA2I1X1 g92565(.B (n_6137), .AN (alu_2nd_operand[9]), .Q (n_302));
  OR2X1 g92566(.A (alu_2nd_operand[10]), .B (n_228), .Q (n_301));
  INX1 g92567(.A (n_290), .Q (n_300));
  NO2X1 g92568(.A (alu_2nd_operand[7]), .B (n_227), .Q (n_299));
  NO2X1 g92569(.A (alu_2nd_operand[6]), .B (n_434), .Q (n_298));
  AN222X1 g49785(.A (alu_2nd_operand[6]), .B (n_434), .C (n_330), .D
       (alu_2nd_operand[5]), .E (n_333), .F (n_226), .Q (n_297));
  AN221X1 g92570(.A (n_233), .B (alu_2nd_operand[8]), .C (n_227), .D
       (alu_2nd_operand[7]), .E (n_303), .Q (n_296));
  NA3I1X0 g50538(.B (n_6134), .C (n_944), .AN (n_8301), .Q (n_295));
  NA2I1X1 g92571(.B (alu_2nd_operand[0]), .AN (n_6121), .Q (n_294));
  NO2X1 g92572(.A (alu_2nd_operand[0]), .B (n_6121), .Q (n_293));
  AN222X1 g92573(.A (csr_data_out[0]), .B (n_8157), .C (n_8166), .D
       (n_7692), .E (n_8296), .F (n_7282), .Q (n_292));
  AN221X1 g49870(.A (n_362), .B (n_6139), .C (n_225), .D
       (alu_2nd_operand[10]), .E (n_224), .Q (n_291));
  NO2I1X1 g92574(.B (alu_2nd_operand[11]), .AN (\rs1_data[11]_39506 ),
       .Q (n_290));
  AO222X1 g92575(.A (n_8166), .B (n_7691), .C (n_8157), .D
       (csr_data_out[11]), .E (n_7935), .F (n_2548), .Q (n_289));
  ON21X1 g50329(.A (alu_2nd_operand[12]), .B (n_432), .C (n_430), .Q
       (n_288));
  ON221X1 g50227(.A (n_161), .B (n_450), .C (n_432), .D
       (\rs1_data[12]_39516 ), .E (n_430), .Q (n_287));
  AO222X1 g92576(.A (n_8166), .B (n_7690), .C (n_8157), .D
       (csr_data_out[12]), .E (n_7936), .F (n_2548), .Q (n_286));
  NA2X1 g92577(.A (n_617), .B (read_data[31]), .Q (n_285));
  AN221X1 g49828(.A (n_405), .B (n_451), .C (n_6155), .D (n_223), .E
       (n_222), .Q (n_284));
  ON21X1 g50555(.A (n_844), .B (n_315), .C (n_405), .Q (n_283));
  ON21X1 g50514(.A (n_8495), .B (n_6132), .C (n_362), .Q (n_282));
  AN321X1 g50221(.A (n_361), .B (n_6132), .C (n_8495), .D (n_8157), .E
       (csr_data_out[16]), .F (n_221), .Q (n_281));
  NO2X1 g92578(.A (n_220), .B (n_219), .Q (n_280));
  INX1 g50328(.A (n_436), .Q (n_279));
  NA2X1 g50539(.A (alu_2nd_operand[17]), .B (n_361), .Q (n_278));
  AO222X1 g92579(.A (read_data[17]), .B (n_160), .C (n_8166), .D
       (n_7685), .E (n_7941), .F (n_2548), .Q (n_277));
  ON21X1 g50365(.A (alu_2nd_operand[18]), .B (n_432), .C (n_430), .Q
       (n_276));
  ON221X1 g50228(.A (n_161), .B (n_650), .C (n_432), .D (n_6141), .E
       (n_430), .Q (n_275));
  AO222X1 g92580(.A (read_data[18]), .B (n_160), .C (n_8166), .D
       (n_7684), .E (n_7942), .F (n_2548), .Q (n_274));
  AN221X1 g49859(.A (n_405), .B (n_649), .C (\rs1_data[19]_39596 ), .D
       (n_218), .E (n_217), .Q (n_273));
  NA2X1 g92581(.A (alu_2nd_operand[1]), .B (n_395), .Q (n_272));
  AN222X0 g50898(.A (n_8166), .B (n_7682), .C (program_counter[1]), .D
       (n_2548), .E (csr_data_out[1]), .F (n_8157), .Q (n_271));
  ON21X1 g50556(.A (alu_2nd_operand[1]), .B (n_6167), .C (n_362), .Q
       (n_270));
  NA2X1 g50575(.A (n_819), .B (n_830), .Q (n_269));
  AND3X1 g49865(.A (n_216), .B (n_215), .C (n_214), .Q (n_268));
  ON211X1 g50212(.A (alu_2nd_operand[21]), .B (n_432), .C (n_430), .D
       (n_213), .Q (n_267));
  AO221X1 g50361(.A (n_362), .B (alu_2nd_operand[21]), .C
       (csr_data_out[21]), .D (n_8157), .E (n_212), .Q (n_266));
  AND4X1 g50634(.A (n_748), .B (n_706), .C (n_743), .D (n_502), .Q
       (n_265));
  AND3X1 g49839(.A (n_211), .B (n_210), .C (n_209), .Q (n_264));
  NA2X1 g50547(.A (alu_2nd_operand[23]), .B (n_361), .Q (n_263));
  AN221X1 g50362(.A (n_8157), .B (csr_data_out[23]), .C
       (alu_2nd_operand[23]), .D (n_362), .E (n_208), .Q (n_262));
  AO222X1 g92582(.A (read_data[24]), .B (n_160), .C (n_8166), .D
       (n_7677), .E (n_7948), .F (n_2548), .Q (n_261));
  AND4X1 g50637(.A (n_579), .B (n_619), .C (n_397), .D (n_690), .Q
       (n_260));
  AO222X1 g92583(.A (read_data[25]), .B (n_160), .C (n_8166), .D
       (n_7676), .E (n_7950), .F (n_2548), .Q (n_259));
  OA211X1 g50568(.A (n_207), .B (alu_2nd_operand[1]), .C (n_505), .D
       (n_744), .Q (n_258));
  NO2X1 g50524(.A (alu_2nd_operand[27]), .B (n_432), .Q (n_257));
  AO222X1 g92584(.A (read_data[27]), .B (n_160), .C (n_8166), .D
       (n_7674), .E (n_7952), .F (n_2548), .Q (n_256));
  AND3X1 g49857(.A (n_206), .B (n_205), .C (n_204), .Q (n_255));
  ON221X1 g50172(.A (n_494), .B (n_376), .C (n_462), .D (n_778), .E
       (n_203), .Q (n_254));
  ON211X1 g50211(.A (alu_2nd_operand[29]), .B (n_432), .C (n_202), .D
       (n_430), .Q (n_253));
  AO221X1 g50360(.A (n_362), .B (alu_2nd_operand[29]), .C
       (csr_data_out[29]), .D (n_8157), .E (n_201), .Q (n_252));
  OA211X1 g92585(.A (n_166), .B (n_686), .C (n_242), .D (n_637), .Q
       (n_251));
  ON221X1 g50229(.A (n_161), .B (n_686), .C (n_432), .D
       (\rs1_data[30]_39526 ), .E (n_430), .Q (n_250));
  AO222X1 g92586(.A (read_data[30]), .B (n_160), .C (n_8166), .D
       (n_7671), .E (n_7955), .F (n_2548), .Q (n_249));
  AN31X1 g49918(.A (n_361), .B (n_6134), .C (alu_2nd_operand[31]), .D
       (n_200), .Q (n_246));
  ON21X1 g50563(.A (alu_2nd_operand[31]), .B (n_6134), .C (n_362), .Q
       (n_245));
  NO2X1 g92589(.A (n_173), .B (n_6181), .Q (n_244));
  AO222X1 g92590(.A (n_8157), .B (csr_data_out[3]), .C (n_8166), .D
       (n_7680), .E (n_7926), .F (n_2548), .Q (n_243));
  NA2X1 g92591(.A (n_530), .B (n_6135), .Q (n_242));
  ON221X1 g50233(.A (n_161), .B (n_497), .C (n_432), .D (n_6178), .E
       (n_430), .Q (n_241));
  AO222X1 g92592(.A (n_8157), .B (csr_data_out[4]), .C (n_8166), .D
       (n_2437), .E (n_7927), .F (n_2548), .Q (n_240));
  ON221X1 g50235(.A (n_161), .B (n_330), .C (n_432), .D (n_6170), .E
       (n_430), .Q (n_239));
  AO222X1 g92593(.A (n_8166), .B (n_8257), .C (n_8157), .D
       (csr_data_out[5]), .E (n_7929), .F (n_2548), .Q (n_238));
  ON221X1 g50231(.A (n_161), .B (n_434), .C (n_432), .D (n_6165), .E
       (n_430), .Q (n_237));
  AO222X1 g92594(.A (n_8166), .B (n_8258), .C (n_8157), .D
       (csr_data_out[6]), .E (n_7930), .F (n_2548), .Q (n_236));
  ON221X1 g50232(.A (n_161), .B (n_227), .C (n_432), .D (n_6183), .E
       (n_430), .Q (n_235));
  AO222X1 g92595(.A (n_8166), .B (n_8259), .C (n_8157), .D
       (csr_data_out[7]), .E (n_7931), .F (n_2548), .Q (n_234));
  INX1 g92596(.A (n_6127), .Q (n_233));
  ON221X0 g50234(.A (n_161), .B (n_233), .C (n_432), .D (n_6127), .E
       (n_430), .Q (n_232));
  AO222X1 g92597(.A (n_8166), .B (n_8260), .C (n_8157), .D
       (csr_data_out[8]), .E (n_7932), .F (n_2548), .Q (n_231));
  AO222X1 g92598(.A (n_8166), .B (n_8261), .C (n_8157), .D
       (csr_data_out[9]), .E (n_7933), .F (n_2548), .Q (n_230));
  INX1 g92599(.A (n_6132), .Q (n_229));
  INX1 g51931(.A (n_6139), .Q (n_228));
  INX1 g92600(.A (n_6183), .Q (n_227));
  ON21X1 g49845(.A (n_831), .B (n_6178), .C (n_199), .Q (n_226));
  ON221X1 g50230(.A (n_161), .B (n_228), .C (n_432), .D (n_6139), .E
       (n_430), .Q (n_225));
  AO222X1 g92601(.A (n_8166), .B (n_8262), .C (n_8157), .D
       (csr_data_out[10]), .E (n_7934), .F (n_2548), .Q (n_224));
  ON221X1 g50208(.A (n_161), .B (n_198), .C (n_432), .D
       (alu_2nd_operand[15]), .E (n_430), .Q (n_223));
  NA3X1 g49916(.A (n_408), .B (n_197), .C (n_196), .Q (n_222));
  AO222X1 g92602(.A (read_data[16]), .B (n_160), .C (n_8166), .D
       (n_7686), .E (n_7940), .F (n_2548), .Q (n_221));
  MU2IX1 g92603(.S (n_8566), .IN0 (read_data[15]), .IN1
       (read_data[31]), .Q (n_220));
  NA2X1 g92604(.A (n_852), .B (n_8162), .Q (n_219));
  ON211X1 g50207(.A (alu_2nd_operand[19]), .B (n_432), .C (n_430), .D
       (n_195), .Q (n_218));
  AO221X1 g50357(.A (n_362), .B (alu_2nd_operand[19]), .C
       (csr_data_out[19]), .D (n_8157), .E (n_194), .Q (n_217));
  ON21X1 g50552(.A (n_472), .B (n_308), .C (n_405), .Q (n_216));
  ON21X1 g50528(.A (alu_2nd_operand[20]), .B (n_6149), .C (n_362), .Q
       (n_215));
  AN321X1 g50214(.A (n_361), .B (n_6149), .C (alu_2nd_operand[20]), .D
       (n_8157), .E (csr_data_out[20]), .F (n_193), .Q (n_214));
  NA2X1 g50549(.A (alu_2nd_operand[21]), .B (n_361), .Q (n_213));
  AO222X1 g92605(.A (read_data[21]), .B (n_160), .C (n_8166), .D
       (n_7693), .E (n_7945), .F (n_2548), .Q (n_212));
  ON21X1 g50550(.A (n_473), .B (n_306), .C (n_405), .Q (n_211));
  ON21X1 g50530(.A (alu_2nd_operand[22]), .B (n_6159), .C (n_362), .Q
       (n_210));
  AN321X1 g50213(.A (n_361), .B (n_6159), .C (alu_2nd_operand[22]), .D
       (n_8157), .E (csr_data_out[22]), .F (n_192), .Q (n_209));
  AO222X1 g92606(.A (read_data[23]), .B (n_160), .C (n_8166), .D
       (n_7678), .E (n_7947), .F (n_2548), .Q (n_208));
  MU2IX1 g92607(.S (alu_2nd_operand[0]), .IN0 (n_6161), .IN1
       (\rs1_data[25]_39346 ), .Q (n_207));
  ON21X1 g50554(.A (n_470), .B (n_309), .C (n_405), .Q (n_206));
  ON21X1 g50526(.A (alu_2nd_operand[28]), .B (n_6136), .C (n_362), .Q
       (n_205));
  AN321X1 g50216(.A (n_361), .B (n_6136), .C (alu_2nd_operand[28]), .D
       (n_8157), .E (csr_data_out[28]), .F (n_191), .Q (n_204));
  OA32X1 g50521(.A (n_498), .B (alu_2nd_operand[0]), .C (n_353), .D
       (n_207), .E (n_780), .Q (n_203));
  NA2X1 g50542(.A (alu_2nd_operand[29]), .B (n_361), .Q (n_202));
  AO222X1 g92608(.A (read_data[29]), .B (n_160), .C (n_8166), .D
       (n_7672), .E (n_7954), .F (n_2548), .Q (n_201));
  NA3X1 g50225(.A (n_436), .B (n_190), .C (n_189), .Q (n_200));
  ON221X1 g49911(.A (n_244), .B (n_188), .C (n_631), .D
       (alu_2nd_operand[3]), .E (n_335), .Q (n_199));
  INX1 g92609(.A (alu_2nd_operand[15]), .Q (n_198));
  NA2X1 g50562(.A (alu_2nd_operand[15]), .B (n_362), .Q (n_197));
  AN222X1 g92610(.A (n_8166), .B (n_7687), .C (n_7939), .D (n_2548), .E
       (csr_data_out[15]), .F (n_8157), .Q (n_196));
  NA2X1 g50561(.A (alu_2nd_operand[19]), .B (n_361), .Q (n_195));
  AO222X1 g92611(.A (read_data[19]), .B (n_160), .C (n_8166), .D
       (n_7683), .E (n_7943), .F (n_2548), .Q (n_194));
  AO222X1 g92612(.A (read_data[20]), .B (n_160), .C (n_8166), .D
       (n_7670), .E (n_7944), .F (n_2548), .Q (n_193));
  AO222X1 g92613(.A (read_data[22]), .B (n_160), .C (n_8166), .D
       (n_7669), .E (n_7946), .F (n_2548), .Q (n_192));
  AO222X1 g92614(.A (read_data[28]), .B (n_160), .C (n_8166), .D
       (n_7673), .E (n_7953), .F (n_2548), .Q (n_191));
  NA2X1 g92615(.A (csr_data_out[31]), .B (n_8157), .Q (n_190));
  AN222X1 g92616(.A (read_data[31]), .B (n_160), .C (n_8166), .D
       (n_8263), .E (n_2548), .F (n_7956), .Q (n_189));
  AN21X1 g50541(.A (n_187), .B (n_347), .C (n_186), .Q (n_188));
  NA2X1 g92617(.A (n_185), .B (n_777), .Q (n_187));
  INX1 g92618(.A (n_348), .Q (n_186));
  NA2X1 g92619(.A (n_272), .B (n_294), .Q (n_185));
  DFRQX1 csr_mcause_interrupt_flag_reg(.C (rc_gclk_199992), .D (n_157),
       .Q (csr_mcause_interrupt_flag));
  DFRQX1 \csr_mcycle_reg[0] (.C (clock), .D (n_2227), .Q
       (csr_mcycle[0]));
  DFRQX1 \csr_mcycle_reg[11] (.C (clock), .D (n_2225), .Q
       (csr_mcycle[11]));
  DFRQX1 \csr_mcycle_reg[12] (.C (clock), .D (n_2224), .Q
       (csr_mcycle[12]));
  DFRQX1 \csr_mcycle_reg[13] (.C (clock), .D (n_2223), .Q
       (csr_mcycle[13]));
  DFRQX2 \csr_mcycle_reg[14] (.C (clock), .D (n_2222), .Q
       (csr_mcycle[14]));
  DFRQX1 \csr_mcycle_reg[15] (.C (clock), .D (n_2221), .Q
       (csr_mcycle[15]));
  DFRQX1 \csr_mcycle_reg[19] (.C (clock), .D (n_2217), .Q
       (csr_mcycle[19]));
  DFRQX1 \csr_mcycle_reg[1] (.C (clock), .D (n_2216), .Q
       (csr_mcycle[1]));
  DFRQX1 \csr_mcycle_reg[21] (.C (clock), .D (n_2214), .Q
       (csr_mcycle[21]));
  DFRQX2 \csr_mcycle_reg[22] (.C (clock), .D (n_2213), .Q
       (csr_mcycle[22]));
  DFRQX1 \csr_mcycle_reg[23] (.C (clock), .D (n_2212), .Q
       (csr_mcycle[23]));
  DFRQX1 \csr_mcycle_reg[24] (.C (clock), .D (n_2211), .Q
       (csr_mcycle[24]));
  DFRQX1 \csr_mcycle_reg[25] (.C (clock), .D (n_2210), .Q
       (csr_mcycle[25]));
  DFRQX1 \csr_mcycle_reg[26] (.C (clock), .D (n_2209), .Q
       (csr_mcycle[26]));
  DFRQX1 \csr_mcycle_reg[27] (.C (clock), .D (n_2208), .Q
       (csr_mcycle[27]));
  DFRQX1 \csr_mcycle_reg[28] (.C (clock), .D (n_2207), .Q
       (csr_mcycle[28]));
  DFRQX1 \csr_mcycle_reg[29] (.C (clock), .D (n_2206), .Q
       (csr_mcycle[29]));
  DFRQX2 \csr_mcycle_reg[2] (.C (clock), .D (n_2205), .Q
       (csr_mcycle[2]));
  DFRQX1 \csr_mcycle_reg[31] (.C (clock), .D (n_2203), .Q
       (csr_mcycle[31]));
  DFRQX2 \csr_mcycle_reg[36] (.C (clock), .D (n_2198), .Q
       (csr_mcycle[36]));
  DFRQX1 \csr_mcycle_reg[3] (.C (clock), .D (n_2194), .Q
       (csr_mcycle[3]));
  DFRQX2 \csr_mcycle_reg[48] (.C (clock), .D (n_2185), .Q
       (csr_mcycle[48]));
  DFRQX1 \csr_mcycle_reg[4] (.C (clock), .D (n_2183), .Q
       (csr_mcycle[4]));
  DFRQX2 \csr_mcycle_reg[50] (.C (clock), .D (n_2182), .Q
       (csr_mcycle[50]));
  DFRQX2 \csr_mcycle_reg[53] (.C (clock), .D (n_2179), .Q
       (csr_mcycle[53]));
  DFRQX2 \csr_mcycle_reg[54] (.C (clock), .D (n_2178), .Q
       (csr_mcycle[54]));
  DFRQX2 \csr_mcycle_reg[56] (.C (clock), .D (n_2176), .Q
       (csr_mcycle[56]));
  DFRQX2 \csr_mcycle_reg[58] (.C (clock), .D (n_2174), .Q
       (csr_mcycle[58]));
  DFRQX1 \csr_mcycle_reg[5] (.C (clock), .D (n_2172), .Q
       (csr_mcycle[5]));
  DFRQX2 \csr_mcycle_reg[60] (.C (clock), .D (n_2171), .Q
       (csr_mcycle[60]));
  DFRQX2 \csr_mcycle_reg[61] (.C (clock), .D (n_2170), .Q
       (csr_mcycle[61]));
  DFRQX2 \csr_mcycle_reg[63] (.C (clock), .D (n_2168), .Q
       (csr_mcycle[63]));
  DFRQX1 \csr_mcycle_reg[7] (.C (clock), .D (n_2166), .Q
       (csr_mcycle[7]));
  DFRQX1 \csr_mcycle_reg[9] (.C (clock), .D (n_2164), .Q
       (csr_mcycle[9]));
  DFRQX1 \csr_mepc_reg[10] (.C (rc_gclk_199945), .D (n_2163), .Q
       (n_7897));
  DFRQX1 \csr_mepc_reg[11] (.C (rc_gclk_199945), .D (n_2162), .Q
       (n_7898));
  DFRQX1 \csr_mepc_reg[12] (.C (rc_gclk_199945), .D (n_2161), .Q
       (n_7899));
  DFRQX1 \csr_mepc_reg[13] (.C (rc_gclk_199945), .D (n_2160), .Q
       (n_7901));
  DFRQX1 \csr_mepc_reg[14] (.C (rc_gclk_199945), .D (n_2159), .Q
       (n_7902));
  DFRQX1 \csr_mepc_reg[15] (.C (rc_gclk_199945), .D (n_2158), .Q
       (n_7903));
  DFRQX1 \csr_mepc_reg[16] (.C (rc_gclk_199945), .D (n_2157), .Q
       (n_7904));
  DFRQX1 \csr_mepc_reg[17] (.C (rc_gclk_199945), .D (n_2156), .Q
       (n_7905));
  DFRQX1 \csr_mepc_reg[18] (.C (rc_gclk_199945), .D (n_2155), .Q
       (n_7906));
  DFRQX1 \csr_mepc_reg[19] (.C (rc_gclk_199945), .D (n_2154), .Q
       (n_7907));
  DFRQX1 \csr_mepc_reg[20] (.C (rc_gclk_199945), .D (n_2153), .Q
       (n_7908));
  DFRQX1 \csr_mepc_reg[21] (.C (rc_gclk_199945), .D (n_2152), .Q
       (n_7909));
  DFRQX1 \csr_mepc_reg[22] (.C (rc_gclk_199945), .D (n_2151), .Q
       (n_7910));
  DFRQX1 \csr_mepc_reg[23] (.C (rc_gclk_199945), .D (n_2150), .Q
       (n_7884));
  DFRQX1 \csr_mepc_reg[24] (.C (rc_gclk_199945), .D (n_2149), .Q
       (n_7885));
  DFRQX1 \csr_mepc_reg[25] (.C (rc_gclk_199945), .D (n_2148), .Q
       (n_7886));
  DFRQX1 \csr_mepc_reg[26] (.C (rc_gclk_199945), .D (n_2147), .Q
       (n_7887));
  DFRQX1 \csr_mepc_reg[27] (.C (rc_gclk_199945), .D (n_2146), .Q
       (n_7888));
  DFRQX1 \csr_mepc_reg[28] (.C (rc_gclk_199945), .D (n_2145), .Q
       (n_7889));
  DFRQX1 \csr_mepc_reg[29] (.C (rc_gclk_199945), .D (n_2144), .Q
       (n_7891));
  DFRQX1 \csr_mepc_reg[2] (.C (rc_gclk_199945), .D (n_2143), .Q
       (n_7890));
  DFRQX1 \csr_mepc_reg[30] (.C (rc_gclk_199945), .D (n_2142), .Q
       (n_7900));
  DFRQX1 \csr_mepc_reg[31] (.C (rc_gclk_199945), .D (n_2141), .Q
       (n_7911));
  DFRQX1 \csr_mepc_reg[3] (.C (rc_gclk_199945), .D (n_2140), .Q
       (n_7964));
  DFRQX1 \csr_mepc_reg[4] (.C (rc_gclk_199945), .D (n_2139), .Q
       (n_7892));
  DFRQX1 \csr_mepc_reg[5] (.C (rc_gclk_199945), .D (n_2138), .Q
       (n_7893));
  DFRQX1 \csr_mepc_reg[6] (.C (rc_gclk_199945), .D (n_2137), .Q
       (n_7894));
  DFRQX1 \csr_mepc_reg[7] (.C (rc_gclk_199945), .D (n_2136), .Q
       (n_7923));
  DFRQX1 \csr_mepc_reg[8] (.C (rc_gclk_199945), .D (n_2135), .Q
       (n_7895));
  DFRQX1 \csr_mepc_reg[9] (.C (rc_gclk_199945), .D (n_2134), .Q
       (n_7896));
  DFRQX1 csr_mie_meie_reg(.C (rc_gclk_199990), .D (n_146), .Q (n_8028));
  DFRQX1 \csr_mie_mfie_reg[0] (.C (rc_gclk_199990), .D (n_116), .Q
       (n_8031));
  DFRQX1 \csr_mie_mfie_reg[10] (.C (rc_gclk_199990), .D (n_2133), .Q
       (n_8043));
  DFRQX1 \csr_mie_mfie_reg[11] (.C (rc_gclk_199990), .D (n_130), .Q
       (n_8045));
  DFRQX1 \csr_mie_mfie_reg[12] (.C (rc_gclk_199990), .D (n_129), .Q
       (n_8046));
  DFRQX1 \csr_mie_mfie_reg[13] (.C (rc_gclk_199990), .D (n_121), .Q
       (n_8047));
  DFRQX1 \csr_mie_mfie_reg[14] (.C (rc_gclk_199990), .D (n_123), .Q
       (n_8048));
  DFRQX1 \csr_mie_mfie_reg[15] (.C (rc_gclk_199990), .D (n_122), .Q
       (n_8049));
  DFRQX1 \csr_mie_mfie_reg[1] (.C (rc_gclk_199990), .D (n_117), .Q
       (n_8033));
  DFRQX1 \csr_mie_mfie_reg[2] (.C (rc_gclk_199990), .D (n_2132), .Q
       (n_8034));
  DFRQX1 \csr_mie_mfie_reg[3] (.C (rc_gclk_199990), .D (n_118), .Q
       (n_8035));
  DFRQX1 \csr_mie_mfie_reg[4] (.C (rc_gclk_199990), .D (n_137), .Q
       (n_8036));
  DFRQX1 \csr_mie_mfie_reg[5] (.C (rc_gclk_199990), .D (n_2131), .Q
       (n_8037));
  DFRQX1 \csr_mie_mfie_reg[6] (.C (rc_gclk_199990), .D (n_2130), .Q
       (n_8039));
  DFRQX1 \csr_mie_mfie_reg[7] (.C (rc_gclk_199990), .D (n_119), .Q
       (n_8040));
  DFRQX1 \csr_mie_mfie_reg[8] (.C (rc_gclk_199990), .D (n_2129), .Q
       (n_8041));
  DFRQX1 \csr_mie_mfie_reg[9] (.C (rc_gclk_199990), .D (n_120), .Q
       (n_8042));
  DFRQX1 csr_mie_msie_reg(.C (rc_gclk_199990), .D (n_115), .Q (n_8030));
  DFRQX1 csr_mie_mtie_reg(.C (rc_gclk_199990), .D (n_2128), .Q
       (n_8029));
  DFRQX1 \csr_minstret_reg[0] (.C (rc_gclk), .D (n_2127), .Q
       (csr_minstret[0]));
  DFRQX1 \csr_minstret_reg[11] (.C (rc_gclk), .D (n_2125), .Q
       (csr_minstret[11]));
  DFRQX1 \csr_minstret_reg[12] (.C (rc_gclk), .D (n_2124), .Q
       (csr_minstret[12]));
  DFRQX1 \csr_minstret_reg[13] (.C (rc_gclk), .D (n_2123), .Q
       (csr_minstret[13]));
  DFRQX1 \csr_minstret_reg[14] (.C (rc_gclk), .D (n_2122), .Q
       (csr_minstret[14]));
  DFRQX1 \csr_minstret_reg[15] (.C (rc_gclk), .D (n_2121), .Q
       (csr_minstret[15]));
  DFRQX1 \csr_minstret_reg[19] (.C (rc_gclk), .D (n_2117), .Q
       (csr_minstret[19]));
  DFRQX1 \csr_minstret_reg[1] (.C (rc_gclk), .D (n_2116), .Q
       (csr_minstret[1]));
  DFRQX1 \csr_minstret_reg[21] (.C (rc_gclk), .D (n_2114), .Q
       (csr_minstret[21]));
  DFRQX1 \csr_minstret_reg[22] (.C (rc_gclk), .D (n_2113), .Q
       (csr_minstret[22]));
  DFRQX1 \csr_minstret_reg[23] (.C (rc_gclk), .D (n_2112), .Q
       (csr_minstret[23]));
  DFRQX1 \csr_minstret_reg[24] (.C (rc_gclk), .D (n_2111), .Q
       (csr_minstret[24]));
  DFRQX1 \csr_minstret_reg[25] (.C (rc_gclk), .D (n_2110), .Q
       (csr_minstret[25]));
  DFRQX1 \csr_minstret_reg[26] (.C (rc_gclk), .D (n_2109), .Q
       (csr_minstret[26]));
  DFRQX1 \csr_minstret_reg[27] (.C (rc_gclk), .D (n_2108), .Q
       (csr_minstret[27]));
  DFRQX1 \csr_minstret_reg[28] (.C (rc_gclk), .D (n_2107), .Q
       (csr_minstret[28]));
  DFRQX1 \csr_minstret_reg[29] (.C (rc_gclk), .D (n_2106), .Q
       (csr_minstret[29]));
  DFRQX1 \csr_minstret_reg[30] (.C (rc_gclk), .D (n_2104), .Q
       (csr_minstret[30]));
  DFRQX1 \csr_minstret_reg[31] (.C (rc_gclk), .D (n_2103), .Q
       (csr_minstret[31]));
  DFRQX2 \csr_minstret_reg[33] (.C (rc_gclk), .D (n_2101), .Q
       (csr_minstret[33]));
  DFRQX1 \csr_minstret_reg[35] (.C (rc_gclk), .D (n_2099), .Q
       (csr_minstret[35]));
  DFRQX1 \csr_minstret_reg[3] (.C (rc_gclk), .D (n_2094), .Q
       (csr_minstret[3]));
  DFRQX2 \csr_minstret_reg[49] (.C (rc_gclk), .D (n_2084), .Q
       (csr_minstret[49]));
  DFRQX1 \csr_minstret_reg[4] (.C (rc_gclk), .D (n_2083), .Q
       (csr_minstret[4]));
  DFRQX2 \csr_minstret_reg[50] (.C (rc_gclk), .D (n_2082), .Q
       (csr_minstret[50]));
  DFRQX2 \csr_minstret_reg[51] (.C (rc_gclk), .D (n_2081), .Q
       (csr_minstret[51]));
  DFRQX2 \csr_minstret_reg[52] (.C (rc_gclk), .D (n_2080), .Q
       (csr_minstret[52]));
  DFRQX2 \csr_minstret_reg[54] (.C (rc_gclk), .D (n_2078), .Q
       (csr_minstret[54]));
  DFRQX2 \csr_minstret_reg[56] (.C (rc_gclk), .D (n_2076), .Q
       (csr_minstret[56]));
  DFRQX2 \csr_minstret_reg[58] (.C (rc_gclk), .D (n_2074), .Q
       (csr_minstret[58]));
  DFRQX1 \csr_minstret_reg[5] (.C (rc_gclk), .D (n_2072), .Q
       (csr_minstret[5]));
  DFRQX2 \csr_minstret_reg[60] (.C (rc_gclk), .D (n_2071), .Q
       (csr_minstret[60]));
  DFRQX2 \csr_minstret_reg[61] (.C (rc_gclk), .D (n_2070), .Q
       (csr_minstret[61]));
  DFRQX2 \csr_minstret_reg[62] (.C (rc_gclk), .D (n_2069), .Q
       (csr_minstret[62]));
  DFRQX2 \csr_minstret_reg[63] (.C (rc_gclk), .D (n_2068), .Q
       (csr_minstret[63]));
  DFRQX2 \csr_minstret_reg[6] (.C (rc_gclk), .D (n_2067), .Q
       (csr_minstret[6]));
  DFRQX1 \csr_minstret_reg[7] (.C (rc_gclk), .D (n_2066), .Q
       (csr_minstret[7]));
  DFRQX1 csr_mstatus_mpie_reg(.C (rc_gclk), .D (n_2056), .Q (n_6256));
  DFRQX1 \csr_mtvec_reg[0] (.C (rc_gclk_199987), .D (n_2023), .Q
       (n_8051));
  DFRQX1 \csr_mtvec_reg[10] (.C (rc_gclk_199987), .D (n_147), .Q
       (csr_mtvec[10]));
  DFRQX1 \csr_mtvec_reg[11] (.C (rc_gclk_199987), .D (n_146), .Q
       (csr_mtvec[11]));
  DFRQX1 \csr_mtvec_reg[12] (.C (rc_gclk_199987), .D (n_2022), .Q
       (csr_mtvec[12]));
  DFRQX1 \csr_mtvec_reg[13] (.C (rc_gclk_199987), .D (n_144), .Q
       (csr_mtvec[13]));
  DFRQX1 \csr_mtvec_reg[14] (.C (rc_gclk_199987), .D (n_143), .Q
       (csr_mtvec[14]));
  DFRQX1 \csr_mtvec_reg[15] (.C (rc_gclk_199987), .D (n_2021), .Q
       (csr_mtvec[15]));
  DFRQX1 \csr_mtvec_reg[16] (.C (rc_gclk_199987), .D (n_116), .Q
       (csr_mtvec[16]));
  DFRQX1 \csr_mtvec_reg[17] (.C (rc_gclk_199987), .D (n_117), .Q
       (csr_mtvec[17]));
  DFRQX1 \csr_mtvec_reg[18] (.C (rc_gclk_199987), .D (n_139), .Q
       (csr_mtvec[18]));
  DFRQX1 \csr_mtvec_reg[19] (.C (rc_gclk_199987), .D (n_118), .Q
       (csr_mtvec[19]));
  DFRQX1 \csr_mtvec_reg[20] (.C (rc_gclk_199987), .D (n_137), .Q
       (csr_mtvec[20]));
  DFRQX1 \csr_mtvec_reg[21] (.C (rc_gclk_199987), .D (n_136), .Q
       (csr_mtvec[21]));
  DFRQX1 \csr_mtvec_reg[22] (.C (rc_gclk_199987), .D (n_135), .Q
       (csr_mtvec[22]));
  DFRQX1 \csr_mtvec_reg[23] (.C (rc_gclk_199987), .D (n_119), .Q
       (csr_mtvec[23]));
  DFRQX1 \csr_mtvec_reg[24] (.C (rc_gclk_199987), .D (n_133), .Q
       (csr_mtvec[24]));
  DFRQX1 \csr_mtvec_reg[25] (.C (rc_gclk_199987), .D (n_120), .Q
       (csr_mtvec[25]));
  DFRQX1 \csr_mtvec_reg[26] (.C (rc_gclk_199987), .D (n_131), .Q
       (csr_mtvec[26]));
  DFRQX1 \csr_mtvec_reg[27] (.C (rc_gclk_199987), .D (n_130), .Q
       (csr_mtvec[27]));
  DFRQX1 \csr_mtvec_reg[28] (.C (rc_gclk_199987), .D (n_2020), .Q
       (csr_mtvec[28]));
  DFRQX1 \csr_mtvec_reg[29] (.C (rc_gclk_199987), .D (n_121), .Q
       (csr_mtvec[29]));
  DFRQX1 \csr_mtvec_reg[2] (.C (rc_gclk_199987), .D (n_2019), .Q
       (csr_mtvec[2]));
  DFRQX1 \csr_mtvec_reg[30] (.C (rc_gclk_199987), .D (n_123), .Q
       (csr_mtvec[30]));
  DFRQX1 \csr_mtvec_reg[31] (.C (rc_gclk_199987), .D (n_122), .Q
       (csr_mtvec[31]));
  DFRQX1 \csr_mtvec_reg[3] (.C (rc_gclk_199987), .D (n_115), .Q
       (csr_mtvec[3]));
  DFRQX1 \csr_mtvec_reg[4] (.C (rc_gclk_199987), .D (n_2018), .Q
       (csr_mtvec[4]));
  DFRQX1 \csr_mtvec_reg[5] (.C (rc_gclk_199987), .D (n_2017), .Q
       (csr_mtvec[5]));
  DFRQX1 \csr_mtvec_reg[6] (.C (rc_gclk_199987), .D (n_2016), .Q
       (csr_mtvec[6]));
  DFRQX1 \csr_mtvec_reg[7] (.C (rc_gclk_199987), .D (n_2015), .Q
       (csr_mtvec[7]));
  DFRQX1 \csr_mtvec_reg[8] (.C (rc_gclk_199987), .D (n_125), .Q
       (csr_mtvec[8]));
  DFRQX1 \csr_mtvec_reg[9] (.C (rc_gclk_199987), .D (n_2014), .Q
       (csr_mtvec[9]));
  DFRQX1 \integer_file_reg[10][0] (.C (rc_gclk_199924), .D (n_2010), .Q
       (n_6464));
  DFRQX1 \integer_file_reg[10][10] (.C (rc_gclk_199924), .D (n_69), .Q
       (n_6805));
  DFRQX1 \integer_file_reg[10][11] (.C (rc_gclk_199924), .D (n_113), .Q
       (n_6836));
  DFRQX1 \integer_file_reg[10][12] (.C (rc_gclk_199924), .D (n_2009),
       .Q (n_6867));
  DFRQX1 \integer_file_reg[10][13] (.C (rc_gclk_199924), .D (n_105), .Q
       (n_6929));
  DFRQX1 \integer_file_reg[10][14] (.C (rc_gclk_199924), .D (n_104), .Q
       (n_6960));
  DFRQX1 \integer_file_reg[10][15] (.C (rc_gclk_199924), .D (n_19), .Q
       (n_6991));
  DFRQX1 \integer_file_reg[10][16] (.C (rc_gclk_199924), .D (n_103), .Q
       (n_7022));
  DFRQX1 \integer_file_reg[10][17] (.C (rc_gclk_199924), .D (n_2008),
       .Q (n_7053));
  DFRQX1 \integer_file_reg[10][18] (.C (rc_gclk_199924), .D (n_56), .Q
       (n_7084));
  DFRQX1 \integer_file_reg[10][19] (.C (rc_gclk_199924), .D (n_2007),
       .Q (n_7115));
  DFRQX1 \integer_file_reg[10][1] (.C (rc_gclk_199924), .D (n_55), .Q
       (n_6495));
  DFRQX1 \integer_file_reg[10][20] (.C (rc_gclk_199924), .D (n_2006),
       .Q (n_7146));
  DFRQX1 \integer_file_reg[10][21] (.C (rc_gclk_199924), .D (n_2005),
       .Q (n_7177));
  DFRQX1 \integer_file_reg[10][22] (.C (rc_gclk_199924), .D (n_2004),
       .Q (n_7208));
  DFRQX1 \integer_file_reg[10][23] (.C (rc_gclk_199924), .D (n_2003),
       .Q (n_6278));
  DFRQX1 \integer_file_reg[10][24] (.C (rc_gclk_199924), .D (n_2002),
       .Q (n_6309));
  DFRQX1 \integer_file_reg[10][25] (.C (rc_gclk_199924), .D (n_2001),
       .Q (n_6340));
  DFRQX1 \integer_file_reg[10][26] (.C (rc_gclk_199924), .D (n_2000),
       .Q (n_6371));
  DFRQX1 \integer_file_reg[10][27] (.C (rc_gclk_199924), .D (n_1999),
       .Q (n_6402));
  DFRQX1 \integer_file_reg[10][28] (.C (rc_gclk_199924), .D (n_1998),
       .Q (n_6433));
  DFRQX1 \integer_file_reg[10][29] (.C (rc_gclk_199924), .D (n_1997),
       .Q (n_6557));
  DFRQX1 \integer_file_reg[10][2] (.C (rc_gclk_199924), .D (n_54), .Q
       (n_6526));
  DFRQX1 \integer_file_reg[10][30] (.C (rc_gclk_199924), .D (n_1996),
       .Q (n_6898));
  DFRQX1 \integer_file_reg[10][31] (.C (rc_gclk_199924), .D (n_1995),
       .Q (n_7239));
  DFRQX1 \integer_file_reg[10][3] (.C (rc_gclk_199924), .D (n_53), .Q
       (n_6588));
  DFRQX1 \integer_file_reg[10][4] (.C (rc_gclk_199924), .D (n_50), .Q
       (n_6619));
  DFRQX1 \integer_file_reg[10][5] (.C (rc_gclk_199924), .D (n_47), .Q
       (n_6650));
  DFRQX1 \integer_file_reg[10][6] (.C (rc_gclk_199924), .D (n_46), .Q
       (n_6681));
  DFRQX1 \integer_file_reg[10][7] (.C (rc_gclk_199924), .D (n_102), .Q
       (n_6712));
  DFRQX1 \integer_file_reg[10][8] (.C (rc_gclk_199924), .D (n_101), .Q
       (n_6743));
  DFRQX1 \integer_file_reg[10][9] (.C (rc_gclk_199924), .D (n_100), .Q
       (n_6774));
  DFRQX1 \integer_file_reg[11][0] (.C (rc_gclk_199948), .D (n_1994), .Q
       (n_6463));
  DFRQX1 \integer_file_reg[11][10] (.C (rc_gclk_199948), .D (n_70), .Q
       (n_6804));
  DFRQX1 \integer_file_reg[11][11] (.C (rc_gclk_199948), .D (n_111), .Q
       (n_6835));
  DFRQX1 \integer_file_reg[11][12] (.C (rc_gclk_199948), .D (n_1993),
       .Q (n_6866));
  DFRQX1 \integer_file_reg[11][13] (.C (rc_gclk_199948), .D (n_108), .Q
       (n_6928));
  DFRQX1 \integer_file_reg[11][14] (.C (rc_gclk_199948), .D (n_104), .Q
       (n_6959));
  DFRQX1 \integer_file_reg[11][15] (.C (rc_gclk_199948), .D (n_19), .Q
       (n_6990));
  DFRQX1 \integer_file_reg[11][16] (.C (rc_gclk_199948), .D (n_98), .Q
       (n_7021));
  DFRQX1 \integer_file_reg[11][17] (.C (rc_gclk_199948), .D (n_91), .Q
       (n_7052));
  DFRQX1 \integer_file_reg[11][18] (.C (rc_gclk_199948), .D (n_56), .Q
       (n_7083));
  DFRQX1 \integer_file_reg[11][19] (.C (rc_gclk_199948), .D (n_1992),
       .Q (n_7114));
  DFRQX1 \integer_file_reg[11][1] (.C (rc_gclk_199948), .D (n_55), .Q
       (n_6494));
  DFRQX1 \integer_file_reg[11][20] (.C (rc_gclk_199948), .D (n_1991),
       .Q (n_7145));
  DFRQX1 \integer_file_reg[11][21] (.C (rc_gclk_199948), .D (n_1990),
       .Q (n_7176));
  DFRQX1 \integer_file_reg[11][22] (.C (rc_gclk_199948), .D (n_1989),
       .Q (n_7207));
  DFRQX1 \integer_file_reg[11][23] (.C (rc_gclk_199948), .D (n_1988),
       .Q (n_6277));
  DFRQX1 \integer_file_reg[11][24] (.C (rc_gclk_199948), .D (n_40), .Q
       (n_6308));
  DFRQX1 \integer_file_reg[11][25] (.C (rc_gclk_199948), .D (n_1987),
       .Q (n_6339));
  DFRQX1 \integer_file_reg[11][26] (.C (rc_gclk_199948), .D (n_6), .Q
       (n_6370));
  DFRQX1 \integer_file_reg[11][27] (.C (rc_gclk_199948), .D (n_1986),
       .Q (n_6401));
  DFRQX1 \integer_file_reg[11][28] (.C (rc_gclk_199948), .D (n_1985),
       .Q (n_6432));
  DFRQX1 \integer_file_reg[11][29] (.C (rc_gclk_199948), .D (n_1984),
       .Q (n_6556));
  DFRQX1 \integer_file_reg[11][2] (.C (rc_gclk_199948), .D (n_39), .Q
       (n_6525));
  DFRQX1 \integer_file_reg[11][30] (.C (rc_gclk_199948), .D (n_1983),
       .Q (n_6897));
  DFRQX1 \integer_file_reg[11][31] (.C (rc_gclk_199948), .D (n_1982),
       .Q (n_7238));
  DFRQX1 \integer_file_reg[11][3] (.C (rc_gclk_199948), .D (n_38), .Q
       (n_6587));
  DFRQX1 \integer_file_reg[11][4] (.C (rc_gclk_199948), .D (n_50), .Q
       (n_6618));
  DFRQX1 \integer_file_reg[11][5] (.C (rc_gclk_199948), .D (n_48), .Q
       (n_6649));
  DFRQX1 \integer_file_reg[11][6] (.C (rc_gclk_199948), .D (n_37), .Q
       (n_6680));
  DFRQX1 \integer_file_reg[11][7] (.C (rc_gclk_199948), .D (n_90), .Q
       (n_6711));
  DFRQX1 \integer_file_reg[11][8] (.C (rc_gclk_199948), .D (n_101), .Q
       (n_6742));
  DFRQX1 \integer_file_reg[11][9] (.C (rc_gclk_199948), .D (n_89), .Q
       (n_6773));
  DFRQX1 \integer_file_reg[12][0] (.C (rc_gclk_199957), .D (n_1981), .Q
       (n_6462));
  DFRQX1 \integer_file_reg[12][10] (.C (rc_gclk_199957), .D (n_36), .Q
       (n_6803));
  DFRQX1 \integer_file_reg[12][11] (.C (rc_gclk_199957), .D (n_110), .Q
       (n_6834));
  DFRQX1 \integer_file_reg[12][12] (.C (rc_gclk_199957), .D (n_1980),
       .Q (n_6865));
  DFRQX1 \integer_file_reg[12][13] (.C (rc_gclk_199957), .D (n_83), .Q
       (n_6927));
  DFRQX1 \integer_file_reg[12][14] (.C (rc_gclk_199957), .D (n_104), .Q
       (n_6958));
  DFRQX1 \integer_file_reg[12][15] (.C (rc_gclk_199957), .D (n_18), .Q
       (n_6989));
  DFRQX1 \integer_file_reg[12][16] (.C (rc_gclk_199957), .D (n_103), .Q
       (n_7020));
  DFRQX1 \integer_file_reg[12][17] (.C (rc_gclk_199957), .D (n_1979),
       .Q (n_7051));
  DFRQX1 \integer_file_reg[12][18] (.C (rc_gclk_199957), .D (n_57), .Q
       (n_7082));
  DFRQX1 \integer_file_reg[12][19] (.C (rc_gclk_199957), .D (n_1978),
       .Q (n_7113));
  DFRQX1 \integer_file_reg[12][1] (.C (rc_gclk_199957), .D (n_55), .Q
       (n_6493));
  DFRQX1 \integer_file_reg[12][20] (.C (rc_gclk_199957), .D (n_1977),
       .Q (n_7144));
  DFRQX1 \integer_file_reg[12][21] (.C (rc_gclk_199957), .D (n_1976),
       .Q (n_7175));
  DFRQX1 \integer_file_reg[12][22] (.C (rc_gclk_199957), .D (n_1975),
       .Q (n_7206));
  DFRQX1 \integer_file_reg[12][23] (.C (rc_gclk_199957), .D (n_1974),
       .Q (n_6276));
  DFRQX1 \integer_file_reg[12][24] (.C (rc_gclk_199957), .D (n_1973),
       .Q (n_6307));
  DFRQX1 \integer_file_reg[12][25] (.C (rc_gclk_199957), .D (n_1972),
       .Q (n_6338));
  DFRQX1 \integer_file_reg[12][26] (.C (rc_gclk_199957), .D (n_6), .Q
       (n_6369));
  DFRQX1 \integer_file_reg[12][27] (.C (rc_gclk_199957), .D (n_1971),
       .Q (n_6400));
  DFRQX1 \integer_file_reg[12][28] (.C (rc_gclk_199957), .D (n_1970),
       .Q (n_6431));
  DFRQX1 \integer_file_reg[12][29] (.C (rc_gclk_199957), .D (n_1969),
       .Q (n_6555));
  DFRQX1 \integer_file_reg[12][2] (.C (rc_gclk_199957), .D (n_39), .Q
       (n_6524));
  DFRQX1 \integer_file_reg[12][30] (.C (rc_gclk_199957), .D (n_1968),
       .Q (n_6896));
  DFRQX1 \integer_file_reg[12][31] (.C (rc_gclk_199957), .D (n_1967),
       .Q (n_7237));
  DFRQX1 \integer_file_reg[12][3] (.C (rc_gclk_199957), .D (n_38), .Q
       (n_6586));
  DFRQX1 \integer_file_reg[12][4] (.C (rc_gclk_199957), .D (n_33), .Q
       (n_6617));
  DFRQX1 \integer_file_reg[12][5] (.C (rc_gclk_199957), .D (n_31), .Q
       (n_6648));
  DFRQX1 \integer_file_reg[12][6] (.C (rc_gclk_199957), .D (n_37), .Q
       (n_6679));
  DFRQX1 \integer_file_reg[12][7] (.C (rc_gclk_199957), .D (n_90), .Q
       (n_6710));
  DFRQX1 \integer_file_reg[12][8] (.C (rc_gclk_199957), .D (n_101), .Q
       (n_6741));
  DFRQX1 \integer_file_reg[12][9] (.C (rc_gclk_199957), .D (n_99), .Q
       (n_6772));
  DFRQX1 \integer_file_reg[13][0] (.C (rc_gclk_199969), .D (n_1966), .Q
       (n_6461));
  DFRQX1 \integer_file_reg[13][10] (.C (rc_gclk_199969), .D (n_36), .Q
       (n_6802));
  DFRQX1 \integer_file_reg[13][11] (.C (rc_gclk_199969), .D (n_112), .Q
       (n_6833));
  DFRQX1 \integer_file_reg[13][12] (.C (rc_gclk_199969), .D (n_1965),
       .Q (n_6864));
  DFRQX1 \integer_file_reg[13][13] (.C (rc_gclk_199969), .D (n_85), .Q
       (n_6926));
  DFRQX1 \integer_file_reg[13][14] (.C (rc_gclk_199969), .D (n_104), .Q
       (n_6957));
  DFRQX1 \integer_file_reg[13][15] (.C (rc_gclk_199969), .D (n_18), .Q
       (n_6988));
  DFRQX1 \integer_file_reg[13][16] (.C (rc_gclk_199969), .D (n_103), .Q
       (n_7019));
  DFRQX1 \integer_file_reg[13][17] (.C (rc_gclk_199969), .D (n_1964),
       .Q (n_7050));
  DFRQX1 \integer_file_reg[13][18] (.C (rc_gclk_199969), .D (n_57), .Q
       (n_7081));
  DFRQX1 \integer_file_reg[13][19] (.C (rc_gclk_199969), .D (n_1963),
       .Q (n_7112));
  DFRQX1 \integer_file_reg[13][1] (.C (rc_gclk_199969), .D (n_30), .Q
       (n_6492));
  DFRQX1 \integer_file_reg[13][20] (.C (rc_gclk_199969), .D (n_1962),
       .Q (n_7143));
  DFRQX1 \integer_file_reg[13][21] (.C (rc_gclk_199969), .D (n_1961),
       .Q (n_7174));
  DFRQX1 \integer_file_reg[13][22] (.C (rc_gclk_199969), .D (n_1960),
       .Q (n_7205));
  DFRQX1 \integer_file_reg[13][23] (.C (rc_gclk_199969), .D (n_1959),
       .Q (n_6275));
  DFRQX1 \integer_file_reg[13][24] (.C (rc_gclk_199969), .D (n_1958),
       .Q (n_6306));
  DFRQX1 \integer_file_reg[13][25] (.C (rc_gclk_199969), .D (n_1957),
       .Q (n_6337));
  DFRQX1 \integer_file_reg[13][26] (.C (rc_gclk_199969), .D (n_7), .Q
       (n_6368));
  DFRQX1 \integer_file_reg[13][27] (.C (rc_gclk_199969), .D (n_1956),
       .Q (n_6399));
  DFRQX1 \integer_file_reg[13][28] (.C (rc_gclk_199969), .D (n_1955),
       .Q (n_6430));
  DFRQX1 \integer_file_reg[13][29] (.C (rc_gclk_199969), .D (n_1954),
       .Q (n_6554));
  DFRQX1 \integer_file_reg[13][2] (.C (rc_gclk_199969), .D (n_54), .Q
       (n_6523));
  DFRQX1 \integer_file_reg[13][30] (.C (rc_gclk_199969), .D (n_1953),
       .Q (n_6895));
  DFRQX1 \integer_file_reg[13][31] (.C (rc_gclk_199969), .D (n_1952),
       .Q (n_7236));
  DFRQX1 \integer_file_reg[13][3] (.C (rc_gclk_199969), .D (n_38), .Q
       (n_6585));
  DFRQX1 \integer_file_reg[13][4] (.C (rc_gclk_199969), .D (n_33), .Q
       (n_6616));
  DFRQX1 \integer_file_reg[13][5] (.C (rc_gclk_199969), .D (n_31), .Q
       (n_6647));
  DFRQX1 \integer_file_reg[13][6] (.C (rc_gclk_199969), .D (n_37), .Q
       (n_6678));
  DFRQX1 \integer_file_reg[13][7] (.C (rc_gclk_199969), .D (n_81), .Q
       (n_6709));
  DFRQX1 \integer_file_reg[13][8] (.C (rc_gclk_199969), .D (n_101), .Q
       (n_6740));
  DFRQX1 \integer_file_reg[13][9] (.C (rc_gclk_199969), .D (n_100), .Q
       (n_6771));
  DFRQX1 \integer_file_reg[14][0] (.C (rc_gclk_199978), .D (n_1951), .Q
       (n_6460));
  DFRQX1 \integer_file_reg[14][10] (.C (rc_gclk_199978), .D (n_36), .Q
       (n_6801));
  DFRQX1 \integer_file_reg[14][11] (.C (rc_gclk_199978), .D (n_112), .Q
       (n_6832));
  DFRQX1 \integer_file_reg[14][12] (.C (rc_gclk_199978), .D (n_1950),
       .Q (n_6863));
  DFRQX1 \integer_file_reg[14][13] (.C (rc_gclk_199978), .D (n_86), .Q
       (n_6925));
  DFRQX1 \integer_file_reg[14][14] (.C (rc_gclk_199978), .D (n_104), .Q
       (n_6956));
  DFRQX1 \integer_file_reg[14][15] (.C (rc_gclk_199978), .D (n_19), .Q
       (n_6987));
  DFRQX1 \integer_file_reg[14][16] (.C (rc_gclk_199978), .D (n_98), .Q
       (n_7018));
  DFRQX1 \integer_file_reg[14][17] (.C (rc_gclk_199978), .D (n_92), .Q
       (n_7049));
  DFRQX1 \integer_file_reg[14][18] (.C (rc_gclk_199978), .D (n_58), .Q
       (n_7080));
  DFRQX1 \integer_file_reg[14][19] (.C (rc_gclk_199978), .D (n_1949),
       .Q (n_7111));
  DFRQX1 \integer_file_reg[14][1] (.C (rc_gclk_199978), .D (n_30), .Q
       (n_6491));
  DFRQX1 \integer_file_reg[14][20] (.C (rc_gclk_199978), .D (n_1948),
       .Q (n_7142));
  DFRQX1 \integer_file_reg[14][21] (.C (rc_gclk_199978), .D (n_1947),
       .Q (n_7173));
  DFRQX1 \integer_file_reg[14][22] (.C (rc_gclk_199978), .D (n_1946),
       .Q (n_7204));
  DFRQX1 \integer_file_reg[14][23] (.C (rc_gclk_199978), .D (n_1945),
       .Q (n_6274));
  DFRQX1 \integer_file_reg[14][24] (.C (rc_gclk_199978), .D (n_1944),
       .Q (n_6305));
  DFRQX1 \integer_file_reg[14][25] (.C (rc_gclk_199978), .D (n_1943),
       .Q (n_6336));
  DFRQX1 \integer_file_reg[14][26] (.C (rc_gclk_199978), .D (n_2), .Q
       (n_6367));
  DFRQX1 \integer_file_reg[14][27] (.C (rc_gclk_199978), .D (n_1942),
       .Q (n_6398));
  DFRQX1 \integer_file_reg[14][28] (.C (rc_gclk_199978), .D (n_1941),
       .Q (n_6429));
  DFRQX1 \integer_file_reg[14][29] (.C (rc_gclk_199978), .D (n_1940),
       .Q (n_6553));
  DFRQX1 \integer_file_reg[14][2] (.C (rc_gclk_199978), .D (n_54), .Q
       (n_6522));
  DFRQX1 \integer_file_reg[14][30] (.C (rc_gclk_199978), .D (n_1939),
       .Q (n_6894));
  DFRQX1 \integer_file_reg[14][31] (.C (rc_gclk_199978), .D (n_1938),
       .Q (n_7235));
  DFRQX1 \integer_file_reg[14][3] (.C (rc_gclk_199978), .D (n_38), .Q
       (n_6584));
  DFRQX1 \integer_file_reg[14][4] (.C (rc_gclk_199978), .D (n_29), .Q
       (n_6615));
  DFRQX1 \integer_file_reg[14][5] (.C (rc_gclk_199978), .D (n_32), .Q
       (n_6646));
  DFRQX1 \integer_file_reg[14][6] (.C (rc_gclk_199978), .D (n_27), .Q
       (n_6677));
  DFRQX1 \integer_file_reg[14][7] (.C (rc_gclk_199978), .D (n_81), .Q
       (n_6708));
  DFRQX1 \integer_file_reg[14][8] (.C (rc_gclk_199978), .D (n_80), .Q
       (n_6739));
  DFRQX1 \integer_file_reg[14][9] (.C (rc_gclk_199978), .D (n_99), .Q
       (n_6770));
  DFRQX1 \integer_file_reg[15][0] (.C (rc_gclk_199888), .D (n_1937), .Q
       (n_6459));
  DFRQX1 \integer_file_reg[15][10] (.C (rc_gclk_199888), .D (n_36), .Q
       (n_6800));
  DFRQX1 \integer_file_reg[15][11] (.C (rc_gclk_199888), .D (n_113), .Q
       (n_6831));
  DFRQX1 \integer_file_reg[15][12] (.C (rc_gclk_199888), .D (n_79), .Q
       (n_6862));
  DFRQX1 \integer_file_reg[15][13] (.C (rc_gclk_199888), .D (n_84), .Q
       (n_6924));
  DFRQX1 \integer_file_reg[15][14] (.C (rc_gclk_199888), .D (n_104), .Q
       (n_6955));
  DFRQX1 \integer_file_reg[15][15] (.C (rc_gclk_199888), .D (n_19), .Q
       (n_6986));
  DFRQX1 \integer_file_reg[15][16] (.C (rc_gclk_199888), .D (n_103), .Q
       (n_7017));
  DFRQX1 \integer_file_reg[15][17] (.C (rc_gclk_199888), .D (n_92), .Q
       (n_7048));
  DFRQX1 \integer_file_reg[15][18] (.C (rc_gclk_199888), .D (n_58), .Q
       (n_7079));
  DFRQX1 \integer_file_reg[15][19] (.C (rc_gclk_199888), .D (n_1936),
       .Q (n_7110));
  DFRQX1 \integer_file_reg[15][1] (.C (rc_gclk_199888), .D (n_26), .Q
       (n_6490));
  DFRQX1 \integer_file_reg[15][20] (.C (rc_gclk_199888), .D (n_1935),
       .Q (n_7141));
  DFRQX1 \integer_file_reg[15][21] (.C (rc_gclk_199888), .D (n_1934),
       .Q (n_7172));
  DFRQX1 \integer_file_reg[15][22] (.C (rc_gclk_199888), .D (n_1933),
       .Q (n_7203));
  DFRQX1 \integer_file_reg[15][23] (.C (rc_gclk_199888), .D (n_1932),
       .Q (n_6273));
  DFRQX1 \integer_file_reg[15][24] (.C (rc_gclk_199888), .D (n_1931),
       .Q (n_6304));
  DFRQX1 \integer_file_reg[15][25] (.C (rc_gclk_199888), .D (n_1930),
       .Q (n_6335));
  DFRQX1 \integer_file_reg[15][26] (.C (rc_gclk_199888), .D (n_7), .Q
       (n_6366));
  DFRQX1 \integer_file_reg[15][27] (.C (rc_gclk_199888), .D (n_1929),
       .Q (n_6397));
  DFRQX1 \integer_file_reg[15][28] (.C (rc_gclk_199888), .D (n_1928),
       .Q (n_6428));
  DFRQX1 \integer_file_reg[15][29] (.C (rc_gclk_199888), .D (n_1927),
       .Q (n_6552));
  DFRQX1 \integer_file_reg[15][2] (.C (rc_gclk_199888), .D (n_39), .Q
       (n_6521));
  DFRQX1 \integer_file_reg[15][30] (.C (rc_gclk_199888), .D (n_1926),
       .Q (n_6893));
  DFRQX1 \integer_file_reg[15][31] (.C (rc_gclk_199888), .D (n_1925),
       .Q (n_7234));
  DFRQX1 \integer_file_reg[15][3] (.C (rc_gclk_199888), .D (n_25), .Q
       (n_6583));
  DFRQX1 \integer_file_reg[15][4] (.C (rc_gclk_199888), .D (n_28), .Q
       (n_6614));
  DFRQX1 \integer_file_reg[15][5] (.C (rc_gclk_199888), .D (n_32), .Q
       (n_6645));
  DFRQX1 \integer_file_reg[15][6] (.C (rc_gclk_199888), .D (n_27), .Q
       (n_6676));
  DFRQX1 \integer_file_reg[15][7] (.C (rc_gclk_199888), .D (n_102), .Q
       (n_6707));
  DFRQX1 \integer_file_reg[15][8] (.C (rc_gclk_199888), .D (n_80), .Q
       (n_6738));
  DFRQX1 \integer_file_reg[15][9] (.C (rc_gclk_199888), .D (n_78), .Q
       (n_6769));
  DFRQX1 \integer_file_reg[16][0] (.C (rc_gclk_199897), .D (n_1924), .Q
       (n_6458));
  DFRQX1 \integer_file_reg[16][10] (.C (rc_gclk_199897), .D (n_36), .Q
       (n_6799));
  DFRQX1 \integer_file_reg[16][11] (.C (rc_gclk_199897), .D (n_111), .Q
       (n_6830));
  DFRQX1 \integer_file_reg[16][12] (.C (rc_gclk_199897), .D (n_77), .Q
       (n_6861));
  DFRQX1 \integer_file_reg[16][13] (.C (rc_gclk_199897), .D (n_76), .Q
       (n_6923));
  DFRQX1 \integer_file_reg[16][14] (.C (rc_gclk_199897), .D (n_104), .Q
       (n_6954));
  DFRQX1 \integer_file_reg[16][15] (.C (rc_gclk_199897), .D (n_19), .Q
       (n_6985));
  DFRQX1 \integer_file_reg[16][16] (.C (rc_gclk_199897), .D (n_103), .Q
       (n_7016));
  DFRQX1 \integer_file_reg[16][17] (.C (rc_gclk_199897), .D (n_93), .Q
       (n_7047));
  DFRQX1 \integer_file_reg[16][18] (.C (rc_gclk_199897), .D (n_59), .Q
       (n_7078));
  DFRQX1 \integer_file_reg[16][19] (.C (rc_gclk_199897), .D (n_1923),
       .Q (n_7109));
  DFRQX1 \integer_file_reg[16][1] (.C (rc_gclk_199897), .D (n_26), .Q
       (n_6489));
  DFRQX1 \integer_file_reg[16][20] (.C (rc_gclk_199897), .D (n_1922),
       .Q (n_7140));
  DFRQX1 \integer_file_reg[16][21] (.C (rc_gclk_199897), .D (n_1921),
       .Q (n_7171));
  DFRQX1 \integer_file_reg[16][22] (.C (rc_gclk_199897), .D (n_1920),
       .Q (n_7202));
  DFRQX1 \integer_file_reg[16][23] (.C (rc_gclk_199897), .D (n_1919),
       .Q (n_6272));
  DFRQX1 \integer_file_reg[16][24] (.C (rc_gclk_199897), .D (n_1918),
       .Q (n_6303));
  DFRQX1 \integer_file_reg[16][25] (.C (rc_gclk_199897), .D (n_1917),
       .Q (n_6334));
  DFRQX1 \integer_file_reg[16][26] (.C (rc_gclk_199897), .D (n_8), .Q
       (n_6365));
  DFRQX1 \integer_file_reg[16][27] (.C (rc_gclk_199897), .D (n_1916),
       .Q (n_6396));
  DFRQX1 \integer_file_reg[16][28] (.C (rc_gclk_199897), .D (n_1915),
       .Q (n_6427));
  DFRQX1 \integer_file_reg[16][29] (.C (rc_gclk_199897), .D (n_1914),
       .Q (n_6551));
  DFRQX1 \integer_file_reg[16][2] (.C (rc_gclk_199897), .D (n_39), .Q
       (n_6520));
  DFRQX1 \integer_file_reg[16][30] (.C (rc_gclk_199897), .D (n_1913),
       .Q (n_6892));
  DFRQX1 \integer_file_reg[16][31] (.C (rc_gclk_199897), .D (n_1912),
       .Q (n_7233));
  DFRQX1 \integer_file_reg[16][3] (.C (rc_gclk_199897), .D (n_53), .Q
       (n_6582));
  DFRQX1 \integer_file_reg[16][4] (.C (rc_gclk_199897), .D (n_33), .Q
       (n_6613));
  DFRQX1 \integer_file_reg[16][5] (.C (rc_gclk_199897), .D (n_32), .Q
       (n_6644));
  DFRQX1 \integer_file_reg[16][6] (.C (rc_gclk_199897), .D (n_27), .Q
       (n_6675));
  DFRQX1 \integer_file_reg[16][7] (.C (rc_gclk_199897), .D (n_102), .Q
       (n_6706));
  DFRQX1 \integer_file_reg[16][8] (.C (rc_gclk_199897), .D (n_80), .Q
       (n_6737));
  DFRQX1 \integer_file_reg[16][9] (.C (rc_gclk_199897), .D (n_99), .Q
       (n_6768));
  DFRQX1 \integer_file_reg[17][0] (.C (rc_gclk_199906), .D (n_1911), .Q
       (n_6457));
  DFRQX1 \integer_file_reg[17][10] (.C (rc_gclk_199906), .D (n_36), .Q
       (n_6798));
  DFRQX1 \integer_file_reg[17][11] (.C (rc_gclk_199906), .D (n_110), .Q
       (n_6829));
  DFRQX1 \integer_file_reg[17][12] (.C (rc_gclk_199906), .D (n_1910),
       .Q (n_6860));
  DFRQX1 \integer_file_reg[17][13] (.C (rc_gclk_199906), .D (n_109), .Q
       (n_6922));
  DFRQX1 \integer_file_reg[17][14] (.C (rc_gclk_199906), .D (n_104), .Q
       (n_6953));
  DFRQX1 \integer_file_reg[17][15] (.C (rc_gclk_199906), .D (n_19), .Q
       (n_6984));
  DFRQX1 \integer_file_reg[17][16] (.C (rc_gclk_199906), .D (n_103), .Q
       (n_7015));
  DFRQX1 \integer_file_reg[17][17] (.C (rc_gclk_199906), .D (n_1909),
       .Q (n_7046));
  DFRQX1 \integer_file_reg[17][18] (.C (rc_gclk_199906), .D (n_59), .Q
       (n_7077));
  DFRQX1 \integer_file_reg[17][19] (.C (rc_gclk_199906), .D (n_1908),
       .Q (n_7108));
  DFRQX1 \integer_file_reg[17][1] (.C (rc_gclk_199906), .D (n_30), .Q
       (n_6488));
  DFRQX1 \integer_file_reg[17][20] (.C (rc_gclk_199906), .D (n_1907),
       .Q (n_7139));
  DFRQX1 \integer_file_reg[17][21] (.C (rc_gclk_199906), .D (n_1906),
       .Q (n_7170));
  DFRQX1 \integer_file_reg[17][22] (.C (rc_gclk_199906), .D (n_1905),
       .Q (n_7201));
  DFRQX1 \integer_file_reg[17][23] (.C (rc_gclk_199906), .D (n_1904),
       .Q (n_6271));
  DFRQX1 \integer_file_reg[17][24] (.C (rc_gclk_199906), .D (n_1903),
       .Q (n_6302));
  DFRQX1 \integer_file_reg[17][25] (.C (rc_gclk_199906), .D (n_1902),
       .Q (n_6333));
  DFRQX1 \integer_file_reg[17][26] (.C (rc_gclk_199906), .D (n_2), .Q
       (n_6364));
  DFRQX1 \integer_file_reg[17][27] (.C (rc_gclk_199906), .D (n_1901),
       .Q (n_6395));
  DFRQX1 \integer_file_reg[17][28] (.C (rc_gclk_199906), .D (n_1900),
       .Q (n_6426));
  DFRQX1 \integer_file_reg[17][29] (.C (rc_gclk_199906), .D (n_1899),
       .Q (n_6550));
  DFRQX1 \integer_file_reg[17][2] (.C (rc_gclk_199906), .D (n_39), .Q
       (n_6519));
  DFRQX1 \integer_file_reg[17][30] (.C (rc_gclk_199906), .D (n_1898),
       .Q (n_6891));
  DFRQX1 \integer_file_reg[17][31] (.C (rc_gclk_199906), .D (n_1897),
       .Q (n_7232));
  DFRQX1 \integer_file_reg[17][3] (.C (rc_gclk_199906), .D (n_53), .Q
       (n_6581));
  DFRQX1 \integer_file_reg[17][4] (.C (rc_gclk_199906), .D (n_35), .Q
       (n_6612));
  DFRQX1 \integer_file_reg[17][5] (.C (rc_gclk_199906), .D (n_31), .Q
       (n_6643));
  DFRQX1 \integer_file_reg[17][6] (.C (rc_gclk_199906), .D (n_27), .Q
       (n_6674));
  DFRQX1 \integer_file_reg[17][7] (.C (rc_gclk_199906), .D (n_81), .Q
       (n_6705));
  DFRQX1 \integer_file_reg[17][8] (.C (rc_gclk_199906), .D (n_80), .Q
       (n_6736));
  DFRQX1 \integer_file_reg[17][9] (.C (rc_gclk_199906), .D (n_99), .Q
       (n_6767));
  DFRQX1 \integer_file_reg[18][0] (.C (rc_gclk_199915), .D (n_1896), .Q
       (n_6456));
  DFRQX1 \integer_file_reg[18][10] (.C (rc_gclk_199915), .D (n_36), .Q
       (n_6797));
  DFRQX1 \integer_file_reg[18][11] (.C (rc_gclk_199915), .D (n_112), .Q
       (n_6828));
  DFRQX1 \integer_file_reg[18][12] (.C (rc_gclk_199915), .D (n_1895),
       .Q (n_6859));
  DFRQX1 \integer_file_reg[18][13] (.C (rc_gclk_199915), .D (n_105), .Q
       (n_6921));
  DFRQX1 \integer_file_reg[18][14] (.C (rc_gclk_199915), .D (n_104), .Q
       (n_6952));
  DFRQX1 \integer_file_reg[18][15] (.C (rc_gclk_199915), .D (n_18), .Q
       (n_6983));
  DFRQX1 \integer_file_reg[18][16] (.C (rc_gclk_199915), .D (n_75), .Q
       (n_7014));
  DFRQX1 \integer_file_reg[18][17] (.C (rc_gclk_199915), .D (n_93), .Q
       (n_7045));
  DFRQX1 \integer_file_reg[18][18] (.C (rc_gclk_199915), .D (n_60), .Q
       (n_7076));
  DFRQX1 \integer_file_reg[18][19] (.C (rc_gclk_199915), .D (n_1894),
       .Q (n_7107));
  DFRQX1 \integer_file_reg[18][1] (.C (rc_gclk_199915), .D (n_24), .Q
       (n_6487));
  DFRQX1 \integer_file_reg[18][20] (.C (rc_gclk_199915), .D (n_1893),
       .Q (n_7138));
  DFRQX1 \integer_file_reg[18][21] (.C (rc_gclk_199915), .D (n_1892),
       .Q (n_7169));
  DFRQX1 \integer_file_reg[18][22] (.C (rc_gclk_199915), .D (n_1891),
       .Q (n_7200));
  DFRQX1 \integer_file_reg[18][23] (.C (rc_gclk_199915), .D (n_1890),
       .Q (n_6270));
  DFRQX1 \integer_file_reg[18][24] (.C (rc_gclk_199915), .D (n_40), .Q
       (n_6301));
  DFRQX1 \integer_file_reg[18][25] (.C (rc_gclk_199915), .D (n_1889),
       .Q (n_6332));
  DFRQX1 \integer_file_reg[18][26] (.C (rc_gclk_199915), .D (n_8), .Q
       (n_6363));
  DFRQX1 \integer_file_reg[18][27] (.C (rc_gclk_199915), .D (n_1888),
       .Q (n_6394));
  DFRQX1 \integer_file_reg[18][28] (.C (rc_gclk_199915), .D (n_1887),
       .Q (n_6425));
  DFRQX1 \integer_file_reg[18][29] (.C (rc_gclk_199915), .D (n_1886),
       .Q (n_6549));
  DFRQX1 \integer_file_reg[18][2] (.C (rc_gclk_199915), .D (n_39), .Q
       (n_6518));
  DFRQX1 \integer_file_reg[18][30] (.C (rc_gclk_199915), .D (n_1885),
       .Q (n_6890));
  DFRQX1 \integer_file_reg[18][31] (.C (rc_gclk_199915), .D (n_1884),
       .Q (n_7231));
  DFRQX1 \integer_file_reg[18][3] (.C (rc_gclk_199915), .D (n_38), .Q
       (n_6580));
  DFRQX1 \integer_file_reg[18][4] (.C (rc_gclk_199915), .D (n_33), .Q
       (n_6611));
  DFRQX1 \integer_file_reg[18][5] (.C (rc_gclk_199915), .D (n_23), .Q
       (n_6642));
  DFRQX1 \integer_file_reg[18][6] (.C (rc_gclk_199915), .D (n_27), .Q
       (n_6673));
  DFRQX1 \integer_file_reg[18][7] (.C (rc_gclk_199915), .D (n_81), .Q
       (n_6704));
  DFRQX1 \integer_file_reg[18][8] (.C (rc_gclk_199915), .D (n_80), .Q
       (n_6735));
  DFRQX1 \integer_file_reg[18][9] (.C (rc_gclk_199915), .D (n_100), .Q
       (n_6766));
  DFRQX1 \integer_file_reg[19][0] (.C (rc_gclk_199927), .D (n_1883), .Q
       (n_6455));
  DFRQX1 \integer_file_reg[19][10] (.C (rc_gclk_199927), .D (n_36), .Q
       (n_6796));
  DFRQX1 \integer_file_reg[19][11] (.C (rc_gclk_199927), .D (n_111), .Q
       (n_6827));
  DFRQX1 \integer_file_reg[19][12] (.C (rc_gclk_199927), .D (n_1882),
       .Q (n_6858));
  DFRQX1 \integer_file_reg[19][13] (.C (rc_gclk_199927), .D (n_85), .Q
       (n_6920));
  DFRQX1 \integer_file_reg[19][14] (.C (rc_gclk_199927), .D (n_104), .Q
       (n_6951));
  DFRQX1 \integer_file_reg[19][15] (.C (rc_gclk_199927), .D (n_18), .Q
       (n_6982));
  DFRQX1 \integer_file_reg[19][16] (.C (rc_gclk_199927), .D (n_75), .Q
       (n_7013));
  DFRQX1 \integer_file_reg[19][17] (.C (rc_gclk_199927), .D (n_94), .Q
       (n_7044));
  DFRQX1 \integer_file_reg[19][18] (.C (rc_gclk_199927), .D (n_60), .Q
       (n_7075));
  DFRQX1 \integer_file_reg[19][19] (.C (rc_gclk_199927), .D (n_1881),
       .Q (n_7106));
  DFRQX1 \integer_file_reg[19][1] (.C (rc_gclk_199927), .D (n_24), .Q
       (n_6486));
  DFRQX1 \integer_file_reg[19][20] (.C (rc_gclk_199927), .D (n_1880),
       .Q (n_7137));
  DFRQX1 \integer_file_reg[19][21] (.C (rc_gclk_199927), .D (n_1879),
       .Q (n_7168));
  DFRQX1 \integer_file_reg[19][22] (.C (rc_gclk_199927), .D (n_1878),
       .Q (n_7199));
  DFRQX1 \integer_file_reg[19][23] (.C (rc_gclk_199927), .D (n_1877),
       .Q (n_6269));
  DFRQX1 \integer_file_reg[19][24] (.C (rc_gclk_199927), .D (n_1876),
       .Q (n_6300));
  DFRQX1 \integer_file_reg[19][25] (.C (rc_gclk_199927), .D (n_1875),
       .Q (n_6331));
  DFRQX1 \integer_file_reg[19][26] (.C (rc_gclk_199927), .D (n_3), .Q
       (n_6362));
  DFRQX1 \integer_file_reg[19][27] (.C (rc_gclk_199927), .D (n_1874),
       .Q (n_6393));
  DFRQX1 \integer_file_reg[19][28] (.C (rc_gclk_199927), .D (n_1873),
       .Q (n_6424));
  DFRQX1 \integer_file_reg[19][29] (.C (rc_gclk_199927), .D (n_1872),
       .Q (n_6548));
  DFRQX1 \integer_file_reg[19][2] (.C (rc_gclk_199927), .D (n_39), .Q
       (n_6517));
  DFRQX1 \integer_file_reg[19][30] (.C (rc_gclk_199927), .D (n_1871),
       .Q (n_6889));
  DFRQX1 \integer_file_reg[19][31] (.C (rc_gclk_199927), .D (n_1870),
       .Q (n_7230));
  DFRQX1 \integer_file_reg[19][3] (.C (rc_gclk_199927), .D (n_38), .Q
       (n_6579));
  DFRQX1 \integer_file_reg[19][4] (.C (rc_gclk_199927), .D (n_29), .Q
       (n_6610));
  DFRQX1 \integer_file_reg[19][5] (.C (rc_gclk_199927), .D (n_23), .Q
       (n_6641));
  DFRQX1 \integer_file_reg[19][6] (.C (rc_gclk_199927), .D (n_27), .Q
       (n_6672));
  DFRQX1 \integer_file_reg[19][7] (.C (rc_gclk_199927), .D (n_82), .Q
       (n_6703));
  DFRQX1 \integer_file_reg[19][8] (.C (rc_gclk_199927), .D (n_80), .Q
       (n_6734));
  DFRQX1 \integer_file_reg[19][9] (.C (rc_gclk_199927), .D (n_78), .Q
       (n_6765));
  DFRQX1 \integer_file_reg[1][0] (.C (rc_gclk_199936), .D (n_1869), .Q
       (n_6473));
  DFRQX1 \integer_file_reg[1][10] (.C (rc_gclk_199936), .D (n_69), .Q
       (n_6814));
  DFRQX1 \integer_file_reg[1][11] (.C (rc_gclk_199936), .D (n_113), .Q
       (n_6845));
  DFRQX1 \integer_file_reg[1][12] (.C (rc_gclk_199936), .D (n_1868), .Q
       (n_6876));
  DFRQX1 \integer_file_reg[1][13] (.C (rc_gclk_199936), .D (n_87), .Q
       (n_6938));
  DFRQX1 \integer_file_reg[1][14] (.C (rc_gclk_199936), .D (n_104), .Q
       (n_6969));
  DFRQX1 \integer_file_reg[1][15] (.C (rc_gclk_199936), .D (n_18), .Q
       (n_7000));
  DFRQX1 \integer_file_reg[1][16] (.C (rc_gclk_199936), .D (n_103), .Q
       (n_7031));
  DFRQX1 \integer_file_reg[1][17] (.C (rc_gclk_199936), .D (n_94), .Q
       (n_7062));
  DFRQX1 \integer_file_reg[1][18] (.C (rc_gclk_199936), .D (n_22), .Q
       (n_7093));
  DFRQX1 \integer_file_reg[1][19] (.C (rc_gclk_199936), .D (n_1867), .Q
       (n_7124));
  DFRQX1 \integer_file_reg[1][1] (.C (rc_gclk_199936), .D (n_30), .Q
       (n_6504));
  DFRQX1 \integer_file_reg[1][20] (.C (rc_gclk_199936), .D (n_1866), .Q
       (n_7155));
  DFRQX1 \integer_file_reg[1][21] (.C (rc_gclk_199936), .D (n_1865), .Q
       (n_7186));
  DFRQX1 \integer_file_reg[1][22] (.C (rc_gclk_199936), .D (n_1864), .Q
       (n_7217));
  DFRQX1 \integer_file_reg[1][23] (.C (rc_gclk_199936), .D (n_1863), .Q
       (n_6287));
  DFRQX1 \integer_file_reg[1][24] (.C (rc_gclk_199936), .D (n_1862), .Q
       (n_6318));
  DFRQX1 \integer_file_reg[1][25] (.C (rc_gclk_199936), .D (n_1861), .Q
       (n_6349));
  DFRQX1 \integer_file_reg[1][26] (.C (rc_gclk_199936), .D (n_9), .Q
       (n_6380));
  DFRQX1 \integer_file_reg[1][27] (.C (rc_gclk_199936), .D (n_1860), .Q
       (n_6411));
  DFRQX1 \integer_file_reg[1][28] (.C (rc_gclk_199936), .D (n_1859), .Q
       (n_6442));
  DFRQX1 \integer_file_reg[1][29] (.C (rc_gclk_199936), .D (n_1858), .Q
       (n_6566));
  DFRQX1 \integer_file_reg[1][2] (.C (rc_gclk_199936), .D (n_39), .Q
       (n_6535));
  DFRQX1 \integer_file_reg[1][30] (.C (rc_gclk_199936), .D (n_1857), .Q
       (n_6907));
  DFRQX1 \integer_file_reg[1][31] (.C (rc_gclk_199936), .D (n_1856), .Q
       (n_7248));
  DFRQX1 \integer_file_reg[1][3] (.C (rc_gclk_199936), .D (n_38), .Q
       (n_6597));
  DFRQX1 \integer_file_reg[1][4] (.C (rc_gclk_199936), .D (n_28), .Q
       (n_6628));
  DFRQX1 \integer_file_reg[1][5] (.C (rc_gclk_199936), .D (n_31), .Q
       (n_6659));
  DFRQX1 \integer_file_reg[1][6] (.C (rc_gclk_199936), .D (n_27), .Q
       (n_6690));
  DFRQX1 \integer_file_reg[1][7] (.C (rc_gclk_199936), .D (n_82), .Q
       (n_6721));
  DFRQX1 \integer_file_reg[1][8] (.C (rc_gclk_199936), .D (n_101), .Q
       (n_6752));
  DFRQX1 \integer_file_reg[1][9] (.C (rc_gclk_199936), .D (n_99), .Q
       (n_6783));
  DFRQX1 \integer_file_reg[20][0] (.C (rc_gclk_199939), .D (n_1855), .Q
       (n_6454));
  DFRQX1 \integer_file_reg[20][10] (.C (rc_gclk_199939), .D (n_70), .Q
       (n_6795));
  DFRQX1 \integer_file_reg[20][11] (.C (rc_gclk_199939), .D (n_111), .Q
       (n_6826));
  DFRQX1 \integer_file_reg[20][12] (.C (rc_gclk_199939), .D (n_79), .Q
       (n_6857));
  DFRQX1 \integer_file_reg[20][13] (.C (rc_gclk_199939), .D (n_106), .Q
       (n_6919));
  DFRQX1 \integer_file_reg[20][14] (.C (rc_gclk_199939), .D (n_104), .Q
       (n_6950));
  DFRQX1 \integer_file_reg[20][15] (.C (rc_gclk_199939), .D (n_18), .Q
       (n_6981));
  DFRQX1 \integer_file_reg[20][16] (.C (rc_gclk_199939), .D (n_103), .Q
       (n_7012));
  DFRQX1 \integer_file_reg[20][17] (.C (rc_gclk_199939), .D (n_95), .Q
       (n_7043));
  DFRQX1 \integer_file_reg[20][18] (.C (rc_gclk_199939), .D (n_22), .Q
       (n_7074));
  DFRQX1 \integer_file_reg[20][19] (.C (rc_gclk_199939), .D (n_1854),
       .Q (n_7105));
  DFRQX1 \integer_file_reg[20][1] (.C (rc_gclk_199939), .D (n_24), .Q
       (n_6485));
  DFRQX1 \integer_file_reg[20][20] (.C (rc_gclk_199939), .D (n_1853),
       .Q (n_7136));
  DFRQX1 \integer_file_reg[20][21] (.C (rc_gclk_199939), .D (n_1852),
       .Q (n_7167));
  DFRQX1 \integer_file_reg[20][22] (.C (rc_gclk_199939), .D (n_1851),
       .Q (n_7198));
  DFRQX1 \integer_file_reg[20][23] (.C (rc_gclk_199939), .D (n_1850),
       .Q (n_6268));
  DFRQX1 \integer_file_reg[20][24] (.C (rc_gclk_199939), .D (n_41), .Q
       (n_6299));
  DFRQX1 \integer_file_reg[20][25] (.C (rc_gclk_199939), .D (n_1849),
       .Q (n_6330));
  DFRQX1 \integer_file_reg[20][26] (.C (rc_gclk_199939), .D (n_9), .Q
       (n_6361));
  DFRQX1 \integer_file_reg[20][27] (.C (rc_gclk_199939), .D (n_1848),
       .Q (n_6392));
  DFRQX1 \integer_file_reg[20][28] (.C (rc_gclk_199939), .D (n_1847),
       .Q (n_6423));
  DFRQX1 \integer_file_reg[20][29] (.C (rc_gclk_199939), .D (n_1846),
       .Q (n_6547));
  DFRQX1 \integer_file_reg[20][2] (.C (rc_gclk_199939), .D (n_21), .Q
       (n_6516));
  DFRQX1 \integer_file_reg[20][30] (.C (rc_gclk_199939), .D (n_1845),
       .Q (n_6888));
  DFRQX1 \integer_file_reg[20][31] (.C (rc_gclk_199939), .D (n_1844),
       .Q (n_7229));
  DFRQX1 \integer_file_reg[20][3] (.C (rc_gclk_199939), .D (n_25), .Q
       (n_6578));
  DFRQX1 \integer_file_reg[20][4] (.C (rc_gclk_199939), .D (n_28), .Q
       (n_6609));
  DFRQX1 \integer_file_reg[20][5] (.C (rc_gclk_199939), .D (n_32), .Q
       (n_6640));
  DFRQX1 \integer_file_reg[20][6] (.C (rc_gclk_199939), .D (n_27), .Q
       (n_6671));
  DFRQX1 \integer_file_reg[20][7] (.C (rc_gclk_199939), .D (n_74), .Q
       (n_6702));
  DFRQX1 \integer_file_reg[20][8] (.C (rc_gclk_199939), .D (n_101), .Q
       (n_6733));
  DFRQX1 \integer_file_reg[20][9] (.C (rc_gclk_199939), .D (n_89), .Q
       (n_6764));
  DFRQX1 \integer_file_reg[21][0] (.C (rc_gclk_199942), .D (n_1843), .Q
       (n_6453));
  DFRQX1 \integer_file_reg[21][10] (.C (rc_gclk_199942), .D (n_70), .Q
       (n_6794));
  DFRQX1 \integer_file_reg[21][11] (.C (rc_gclk_199942), .D (n_110), .Q
       (n_6825));
  DFRQX1 \integer_file_reg[21][12] (.C (rc_gclk_199942), .D (n_79), .Q
       (n_6856));
  DFRQX1 \integer_file_reg[21][13] (.C (rc_gclk_199942), .D (n_108), .Q
       (n_6918));
  DFRQX1 \integer_file_reg[21][14] (.C (rc_gclk_199942), .D (n_73), .Q
       (n_6949));
  DFRQX1 \integer_file_reg[21][15] (.C (rc_gclk_199942), .D (n_18), .Q
       (n_6980));
  DFRQX1 \integer_file_reg[21][16] (.C (rc_gclk_199942), .D (n_75), .Q
       (n_7011));
  DFRQX1 \integer_file_reg[21][17] (.C (rc_gclk_199942), .D (n_95), .Q
       (n_7042));
  DFRQX1 \integer_file_reg[21][18] (.C (rc_gclk_199942), .D (n_61), .Q
       (n_7073));
  DFRQX1 \integer_file_reg[21][19] (.C (rc_gclk_199942), .D (n_1842),
       .Q (n_7104));
  DFRQX1 \integer_file_reg[21][1] (.C (rc_gclk_199942), .D (n_24), .Q
       (n_6484));
  DFRQX1 \integer_file_reg[21][20] (.C (rc_gclk_199942), .D (n_1841),
       .Q (n_7135));
  DFRQX1 \integer_file_reg[21][21] (.C (rc_gclk_199942), .D (n_1840),
       .Q (n_7166));
  DFRQX1 \integer_file_reg[21][22] (.C (rc_gclk_199942), .D (n_1839),
       .Q (n_7197));
  DFRQX1 \integer_file_reg[21][23] (.C (rc_gclk_199942), .D (n_1838),
       .Q (n_6267));
  DFRQX1 \integer_file_reg[21][24] (.C (rc_gclk_199942), .D (n_1837),
       .Q (n_6298));
  DFRQX1 \integer_file_reg[21][25] (.C (rc_gclk_199942), .D (n_1836),
       .Q (n_6329));
  DFRQX1 \integer_file_reg[21][26] (.C (rc_gclk_199942), .D (n_10), .Q
       (n_6360));
  DFRQX1 \integer_file_reg[21][27] (.C (rc_gclk_199942), .D (n_1835),
       .Q (n_6391));
  DFRQX1 \integer_file_reg[21][28] (.C (rc_gclk_199942), .D (n_1834),
       .Q (n_6422));
  DFRQX1 \integer_file_reg[21][29] (.C (rc_gclk_199942), .D (n_1833),
       .Q (n_6546));
  DFRQX1 \integer_file_reg[21][2] (.C (rc_gclk_199942), .D (n_21), .Q
       (n_6515));
  DFRQX1 \integer_file_reg[21][30] (.C (rc_gclk_199942), .D (n_1832),
       .Q (n_6887));
  DFRQX1 \integer_file_reg[21][31] (.C (rc_gclk_199942), .D (n_1831),
       .Q (n_7228));
  DFRQX1 \integer_file_reg[21][3] (.C (rc_gclk_199942), .D (n_25), .Q
       (n_6577));
  DFRQX1 \integer_file_reg[21][4] (.C (rc_gclk_199942), .D (n_29), .Q
       (n_6608));
  DFRQX1 \integer_file_reg[21][5] (.C (rc_gclk_199942), .D (n_32), .Q
       (n_6639));
  DFRQX1 \integer_file_reg[21][6] (.C (rc_gclk_199942), .D (n_37), .Q
       (n_6670));
  DFRQX1 \integer_file_reg[21][7] (.C (rc_gclk_199942), .D (n_74), .Q
       (n_6701));
  DFRQX1 \integer_file_reg[21][8] (.C (rc_gclk_199942), .D (n_80), .Q
       (n_6732));
  DFRQX1 \integer_file_reg[21][9] (.C (rc_gclk_199942), .D (n_78), .Q
       (n_6763));
  DFRQX1 \integer_file_reg[22][0] (.C (rc_gclk_199951), .D (n_1830), .Q
       (n_6452));
  DFRQX1 \integer_file_reg[22][10] (.C (rc_gclk_199951), .D (n_69), .Q
       (n_6793));
  DFRQX1 \integer_file_reg[22][11] (.C (rc_gclk_199951), .D (n_111), .Q
       (n_6824));
  DFRQX1 \integer_file_reg[22][12] (.C (rc_gclk_199951), .D (n_1829),
       .Q (n_6855));
  DFRQX1 \integer_file_reg[22][13] (.C (rc_gclk_199951), .D (n_86), .Q
       (n_6917));
  DFRQX1 \integer_file_reg[22][14] (.C (rc_gclk_199951), .D (n_73), .Q
       (n_6948));
  DFRQX1 \integer_file_reg[22][15] (.C (rc_gclk_199951), .D (n_18), .Q
       (n_6979));
  DFRQX1 \integer_file_reg[22][16] (.C (rc_gclk_199951), .D (n_98), .Q
       (n_7010));
  DFRQX1 \integer_file_reg[22][17] (.C (rc_gclk_199951), .D (n_1828),
       .Q (n_7041));
  DFRQX1 \integer_file_reg[22][18] (.C (rc_gclk_199951), .D (n_22), .Q
       (n_7072));
  DFRQX1 \integer_file_reg[22][19] (.C (rc_gclk_199951), .D (n_1827),
       .Q (n_7103));
  DFRQX1 \integer_file_reg[22][1] (.C (rc_gclk_199951), .D (n_30), .Q
       (n_6483));
  DFRQX1 \integer_file_reg[22][20] (.C (rc_gclk_199951), .D (n_1826),
       .Q (n_7134));
  DFRQX1 \integer_file_reg[22][21] (.C (rc_gclk_199951), .D (n_1825),
       .Q (n_7165));
  DFRQX1 \integer_file_reg[22][22] (.C (rc_gclk_199951), .D (n_1824),
       .Q (n_7196));
  DFRQX1 \integer_file_reg[22][23] (.C (rc_gclk_199951), .D (n_1823),
       .Q (n_6266));
  DFRQX1 \integer_file_reg[22][24] (.C (rc_gclk_199951), .D (n_41), .Q
       (n_6297));
  DFRQX1 \integer_file_reg[22][25] (.C (rc_gclk_199951), .D (n_1822),
       .Q (n_6328));
  DFRQX1 \integer_file_reg[22][26] (.C (rc_gclk_199951), .D (n_10), .Q
       (n_6359));
  DFRQX1 \integer_file_reg[22][27] (.C (rc_gclk_199951), .D (n_1821),
       .Q (n_6390));
  DFRQX1 \integer_file_reg[22][28] (.C (rc_gclk_199951), .D (n_1820),
       .Q (n_6421));
  DFRQX1 \integer_file_reg[22][29] (.C (rc_gclk_199951), .D (n_1819),
       .Q (n_6545));
  DFRQX1 \integer_file_reg[22][2] (.C (rc_gclk_199951), .D (n_39), .Q
       (n_6514));
  DFRQX1 \integer_file_reg[22][30] (.C (rc_gclk_199951), .D (n_1818),
       .Q (n_6886));
  DFRQX1 \integer_file_reg[22][31] (.C (rc_gclk_199951), .D (n_1817),
       .Q (n_7227));
  DFRQX1 \integer_file_reg[22][3] (.C (rc_gclk_199951), .D (n_38), .Q
       (n_6576));
  DFRQX1 \integer_file_reg[22][4] (.C (rc_gclk_199951), .D (n_34), .Q
       (n_6607));
  DFRQX1 \integer_file_reg[22][5] (.C (rc_gclk_199951), .D (n_31), .Q
       (n_6638));
  DFRQX1 \integer_file_reg[22][6] (.C (rc_gclk_199951), .D (n_37), .Q
       (n_6669));
  DFRQX1 \integer_file_reg[22][7] (.C (rc_gclk_199951), .D (n_74), .Q
       (n_6700));
  DFRQX1 \integer_file_reg[22][8] (.C (rc_gclk_199951), .D (n_80), .Q
       (n_6731));
  DFRQX1 \integer_file_reg[22][9] (.C (rc_gclk_199951), .D (n_99), .Q
       (n_6762));
  DFRQX1 \integer_file_reg[23][0] (.C (rc_gclk_199954), .D (n_1816), .Q
       (n_6451));
  DFRQX1 \integer_file_reg[23][10] (.C (rc_gclk_199954), .D (n_70), .Q
       (n_6792));
  DFRQX1 \integer_file_reg[23][11] (.C (rc_gclk_199954), .D (n_112), .Q
       (n_6823));
  DFRQX1 \integer_file_reg[23][12] (.C (rc_gclk_199954), .D (n_1815),
       .Q (n_6854));
  DFRQX1 \integer_file_reg[23][13] (.C (rc_gclk_199954), .D (n_88), .Q
       (n_6916));
  DFRQX1 \integer_file_reg[23][14] (.C (rc_gclk_199954), .D (n_104), .Q
       (n_6947));
  DFRQX1 \integer_file_reg[23][15] (.C (rc_gclk_199954), .D (n_19), .Q
       (n_6978));
  DFRQX1 \integer_file_reg[23][16] (.C (rc_gclk_199954), .D (n_75), .Q
       (n_7009));
  DFRQX1 \integer_file_reg[23][17] (.C (rc_gclk_199954), .D (n_96), .Q
       (n_7040));
  DFRQX1 \integer_file_reg[23][18] (.C (rc_gclk_199954), .D (n_61), .Q
       (n_7071));
  DFRQX1 \integer_file_reg[23][19] (.C (rc_gclk_199954), .D (n_1814),
       .Q (n_7102));
  DFRQX1 \integer_file_reg[23][1] (.C (rc_gclk_199954), .D (n_30), .Q
       (n_6482));
  DFRQX1 \integer_file_reg[23][20] (.C (rc_gclk_199954), .D (n_1813),
       .Q (n_7133));
  DFRQX1 \integer_file_reg[23][21] (.C (rc_gclk_199954), .D (n_1812),
       .Q (n_7164));
  DFRQX1 \integer_file_reg[23][22] (.C (rc_gclk_199954), .D (n_1811),
       .Q (n_7195));
  DFRQX1 \integer_file_reg[23][23] (.C (rc_gclk_199954), .D (n_1810),
       .Q (n_6265));
  DFRQX1 \integer_file_reg[23][24] (.C (rc_gclk_199954), .D (n_42), .Q
       (n_6296));
  DFRQX1 \integer_file_reg[23][25] (.C (rc_gclk_199954), .D (n_1809),
       .Q (n_6327));
  DFRQX1 \integer_file_reg[23][26] (.C (rc_gclk_199954), .D (n_3), .Q
       (n_6358));
  DFRQX1 \integer_file_reg[23][27] (.C (rc_gclk_199954), .D (n_1808),
       .Q (n_6389));
  DFRQX1 \integer_file_reg[23][28] (.C (rc_gclk_199954), .D (n_1807),
       .Q (n_6420));
  DFRQX1 \integer_file_reg[23][29] (.C (rc_gclk_199954), .D (n_1806),
       .Q (n_6544));
  DFRQX1 \integer_file_reg[23][2] (.C (rc_gclk_199954), .D (n_39), .Q
       (n_6513));
  DFRQX1 \integer_file_reg[23][30] (.C (rc_gclk_199954), .D (n_1805),
       .Q (n_6885));
  DFRQX1 \integer_file_reg[23][31] (.C (rc_gclk_199954), .D (n_1804),
       .Q (n_7226));
  DFRQX1 \integer_file_reg[23][3] (.C (rc_gclk_199954), .D (n_25), .Q
       (n_6575));
  DFRQX1 \integer_file_reg[23][4] (.C (rc_gclk_199954), .D (n_33), .Q
       (n_6606));
  DFRQX1 \integer_file_reg[23][5] (.C (rc_gclk_199954), .D (n_48), .Q
       (n_6637));
  DFRQX1 \integer_file_reg[23][6] (.C (rc_gclk_199954), .D (n_37), .Q
       (n_6668));
  DFRQX1 \integer_file_reg[23][7] (.C (rc_gclk_199954), .D (n_74), .Q
       (n_6699));
  DFRQX1 \integer_file_reg[23][8] (.C (rc_gclk_199954), .D (n_72), .Q
       (n_6730));
  DFRQX1 \integer_file_reg[23][9] (.C (rc_gclk_199954), .D (n_100), .Q
       (n_6761));
  DFRQX1 \integer_file_reg[24][0] (.C (rc_gclk_199960), .D (n_1803), .Q
       (n_6450));
  DFRQX1 \integer_file_reg[24][10] (.C (rc_gclk_199960), .D (n_70), .Q
       (n_6791));
  DFRQX1 \integer_file_reg[24][11] (.C (rc_gclk_199960), .D (n_112), .Q
       (n_6822));
  DFRQX1 \integer_file_reg[24][12] (.C (rc_gclk_199960), .D (n_79), .Q
       (n_6853));
  DFRQX1 \integer_file_reg[24][13] (.C (rc_gclk_199960), .D (n_76), .Q
       (n_6915));
  DFRQX1 \integer_file_reg[24][14] (.C (rc_gclk_199960), .D (n_104), .Q
       (n_6946));
  DFRQX1 \integer_file_reg[24][15] (.C (rc_gclk_199960), .D (n_19), .Q
       (n_6977));
  DFRQX1 \integer_file_reg[24][16] (.C (rc_gclk_199960), .D (n_75), .Q
       (n_7008));
  DFRQX1 \integer_file_reg[24][17] (.C (rc_gclk_199960), .D (n_1802),
       .Q (n_7039));
  DFRQX1 \integer_file_reg[24][18] (.C (rc_gclk_199960), .D (n_62), .Q
       (n_7070));
  DFRQX1 \integer_file_reg[24][19] (.C (rc_gclk_199960), .D (n_1801),
       .Q (n_7101));
  DFRQX1 \integer_file_reg[24][1] (.C (rc_gclk_199960), .D (n_24), .Q
       (n_6481));
  DFRQX1 \integer_file_reg[24][20] (.C (rc_gclk_199960), .D (n_1800),
       .Q (n_7132));
  DFRQX1 \integer_file_reg[24][21] (.C (rc_gclk_199960), .D (n_1799),
       .Q (n_7163));
  DFRQX1 \integer_file_reg[24][22] (.C (rc_gclk_199960), .D (n_1798),
       .Q (n_7194));
  DFRQX1 \integer_file_reg[24][23] (.C (rc_gclk_199960), .D (n_1797),
       .Q (n_6264));
  DFRQX1 \integer_file_reg[24][24] (.C (rc_gclk_199960), .D (n_1796),
       .Q (n_6295));
  DFRQX1 \integer_file_reg[24][25] (.C (rc_gclk_199960), .D (n_1795),
       .Q (n_6326));
  DFRQX1 \integer_file_reg[24][26] (.C (rc_gclk_199960), .D (n_4), .Q
       (n_6357));
  DFRQX1 \integer_file_reg[24][27] (.C (rc_gclk_199960), .D (n_1794),
       .Q (n_6388));
  DFRQX1 \integer_file_reg[24][28] (.C (rc_gclk_199960), .D (n_1793),
       .Q (n_6419));
  DFRQX1 \integer_file_reg[24][29] (.C (rc_gclk_199960), .D (n_1792),
       .Q (n_6543));
  DFRQX1 \integer_file_reg[24][2] (.C (rc_gclk_199960), .D (n_54), .Q
       (n_6512));
  DFRQX1 \integer_file_reg[24][30] (.C (rc_gclk_199960), .D (n_1791),
       .Q (n_6884));
  DFRQX1 \integer_file_reg[24][31] (.C (rc_gclk_199960), .D (n_1790),
       .Q (n_7225));
  DFRQX1 \integer_file_reg[24][3] (.C (rc_gclk_199960), .D (n_25), .Q
       (n_6574));
  DFRQX1 \integer_file_reg[24][4] (.C (rc_gclk_199960), .D (n_33), .Q
       (n_6605));
  DFRQX1 \integer_file_reg[24][5] (.C (rc_gclk_199960), .D (n_47), .Q
       (n_6636));
  DFRQX1 \integer_file_reg[24][6] (.C (rc_gclk_199960), .D (n_37), .Q
       (n_6667));
  DFRQX1 \integer_file_reg[24][7] (.C (rc_gclk_199960), .D (n_81), .Q
       (n_6698));
  DFRQX1 \integer_file_reg[24][8] (.C (rc_gclk_199960), .D (n_72), .Q
       (n_6729));
  DFRQX1 \integer_file_reg[24][9] (.C (rc_gclk_199960), .D (n_100), .Q
       (n_6760));
  DFRQX1 \integer_file_reg[25][0] (.C (rc_gclk_199963), .D (n_1789), .Q
       (n_6449));
  DFRQX1 \integer_file_reg[25][10] (.C (rc_gclk_199963), .D (n_70), .Q
       (n_6790));
  DFRQX1 \integer_file_reg[25][11] (.C (rc_gclk_199963), .D (n_111), .Q
       (n_6821));
  DFRQX1 \integer_file_reg[25][12] (.C (rc_gclk_199963), .D (n_77), .Q
       (n_6852));
  DFRQX1 \integer_file_reg[25][13] (.C (rc_gclk_199963), .D (n_87), .Q
       (n_6914));
  DFRQX1 \integer_file_reg[25][14] (.C (rc_gclk_199963), .D (n_71), .Q
       (n_6945));
  DFRQX1 \integer_file_reg[25][15] (.C (rc_gclk_199963), .D (n_18), .Q
       (n_6976));
  DFRQX1 \integer_file_reg[25][16] (.C (rc_gclk_199963), .D (n_98), .Q
       (n_7007));
  DFRQX1 \integer_file_reg[25][17] (.C (rc_gclk_199963), .D (n_96), .Q
       (n_7038));
  DFRQX1 \integer_file_reg[25][18] (.C (rc_gclk_199963), .D (n_62), .Q
       (n_7069));
  DFRQX1 \integer_file_reg[25][19] (.C (rc_gclk_199963), .D (n_1788),
       .Q (n_7100));
  DFRQX1 \integer_file_reg[25][1] (.C (rc_gclk_199963), .D (n_24), .Q
       (n_6480));
  DFRQX1 \integer_file_reg[25][20] (.C (rc_gclk_199963), .D (n_1787),
       .Q (n_7131));
  DFRQX1 \integer_file_reg[25][21] (.C (rc_gclk_199963), .D (n_1786),
       .Q (n_7162));
  DFRQX1 \integer_file_reg[25][22] (.C (rc_gclk_199963), .D (n_1785),
       .Q (n_7193));
  DFRQX1 \integer_file_reg[25][23] (.C (rc_gclk_199963), .D (n_1784),
       .Q (n_6263));
  DFRQX1 \integer_file_reg[25][24] (.C (rc_gclk_199963), .D (n_1783),
       .Q (n_6294));
  DFRQX1 \integer_file_reg[25][25] (.C (rc_gclk_199963), .D (n_1782),
       .Q (n_6325));
  DFRQX1 \integer_file_reg[25][26] (.C (rc_gclk_199963), .D (n_11), .Q
       (n_6356));
  DFRQX1 \integer_file_reg[25][27] (.C (rc_gclk_199963), .D (n_1781),
       .Q (n_6387));
  DFRQX1 \integer_file_reg[25][28] (.C (rc_gclk_199963), .D (n_1780),
       .Q (n_6418));
  DFRQX1 \integer_file_reg[25][29] (.C (rc_gclk_199963), .D (n_1779),
       .Q (n_6542));
  DFRQX1 \integer_file_reg[25][2] (.C (rc_gclk_199963), .D (n_54), .Q
       (n_6511));
  DFRQX1 \integer_file_reg[25][30] (.C (rc_gclk_199963), .D (n_1778),
       .Q (n_6883));
  DFRQX1 \integer_file_reg[25][31] (.C (rc_gclk_199963), .D (n_1777),
       .Q (n_7224));
  DFRQX1 \integer_file_reg[25][3] (.C (rc_gclk_199963), .D (n_25), .Q
       (n_6573));
  DFRQX1 \integer_file_reg[25][4] (.C (rc_gclk_199963), .D (n_52), .Q
       (n_6604));
  DFRQX1 \integer_file_reg[25][5] (.C (rc_gclk_199963), .D (n_31), .Q
       (n_6635));
  DFRQX1 \integer_file_reg[25][6] (.C (rc_gclk_199963), .D (n_46), .Q
       (n_6666));
  DFRQX1 \integer_file_reg[25][7] (.C (rc_gclk_199963), .D (n_81), .Q
       (n_6697));
  DFRQX1 \integer_file_reg[25][8] (.C (rc_gclk_199963), .D (n_80), .Q
       (n_6728));
  DFRQX1 \integer_file_reg[25][9] (.C (rc_gclk_199963), .D (n_89), .Q
       (n_6759));
  DFRQX1 \integer_file_reg[26][0] (.C (rc_gclk_199972), .D (n_1776), .Q
       (n_6448));
  DFRQX1 \integer_file_reg[26][10] (.C (rc_gclk_199972), .D (n_69), .Q
       (n_6789));
  DFRQX1 \integer_file_reg[26][11] (.C (rc_gclk_199972), .D (n_111), .Q
       (n_6820));
  DFRQX1 \integer_file_reg[26][12] (.C (rc_gclk_199972), .D (n_1775),
       .Q (n_6851));
  DFRQX1 \integer_file_reg[26][13] (.C (rc_gclk_199972), .D (n_107), .Q
       (n_6913));
  DFRQX1 \integer_file_reg[26][14] (.C (rc_gclk_199972), .D (n_71), .Q
       (n_6944));
  DFRQX1 \integer_file_reg[26][15] (.C (rc_gclk_199972), .D (n_18), .Q
       (n_6975));
  DFRQX1 \integer_file_reg[26][16] (.C (rc_gclk_199972), .D (n_103), .Q
       (n_7006));
  DFRQX1 \integer_file_reg[26][17] (.C (rc_gclk_199972), .D (n_97), .Q
       (n_7037));
  DFRQX1 \integer_file_reg[26][18] (.C (rc_gclk_199972), .D (n_22), .Q
       (n_7068));
  DFRQX1 \integer_file_reg[26][19] (.C (rc_gclk_199972), .D (n_1774),
       .Q (n_7099));
  DFRQX1 \integer_file_reg[26][1] (.C (rc_gclk_199972), .D (n_30), .Q
       (n_6479));
  DFRQX1 \integer_file_reg[26][20] (.C (rc_gclk_199972), .D (n_1773),
       .Q (n_7130));
  DFRQX1 \integer_file_reg[26][21] (.C (rc_gclk_199972), .D (n_1772),
       .Q (n_7161));
  DFRQX1 \integer_file_reg[26][22] (.C (rc_gclk_199972), .D (n_1771),
       .Q (n_7192));
  DFRQX1 \integer_file_reg[26][23] (.C (rc_gclk_199972), .D (n_1770),
       .Q (n_6262));
  DFRQX1 \integer_file_reg[26][24] (.C (rc_gclk_199972), .D (n_1769),
       .Q (n_6293));
  DFRQX1 \integer_file_reg[26][25] (.C (rc_gclk_199972), .D (n_1768),
       .Q (n_6324));
  DFRQX1 \integer_file_reg[26][26] (.C (rc_gclk_199972), .D (n_11), .Q
       (n_6355));
  DFRQX1 \integer_file_reg[26][27] (.C (rc_gclk_199972), .D (n_1767),
       .Q (n_6386));
  DFRQX1 \integer_file_reg[26][28] (.C (rc_gclk_199972), .D (n_1766),
       .Q (n_6417));
  DFRQX1 \integer_file_reg[26][29] (.C (rc_gclk_199972), .D (n_1765),
       .Q (n_6541));
  DFRQX1 \integer_file_reg[26][2] (.C (rc_gclk_199972), .D (n_39), .Q
       (n_6510));
  DFRQX1 \integer_file_reg[26][30] (.C (rc_gclk_199972), .D (n_1764),
       .Q (n_6882));
  DFRQX1 \integer_file_reg[26][31] (.C (rc_gclk_199972), .D (n_1763),
       .Q (n_7223));
  DFRQX1 \integer_file_reg[26][3] (.C (rc_gclk_199972), .D (n_25), .Q
       (n_6572));
  DFRQX1 \integer_file_reg[26][4] (.C (rc_gclk_199972), .D (n_52), .Q
       (n_6603));
  DFRQX1 \integer_file_reg[26][5] (.C (rc_gclk_199972), .D (n_31), .Q
       (n_6634));
  DFRQX1 \integer_file_reg[26][6] (.C (rc_gclk_199972), .D (n_46), .Q
       (n_6665));
  DFRQX1 \integer_file_reg[26][7] (.C (rc_gclk_199972), .D (n_81), .Q
       (n_6696));
  DFRQX1 \integer_file_reg[26][8] (.C (rc_gclk_199972), .D (n_80), .Q
       (n_6727));
  DFRQX1 \integer_file_reg[26][9] (.C (rc_gclk_199972), .D (n_78), .Q
       (n_6758));
  DFRQX1 \integer_file_reg[27][0] (.C (rc_gclk_199975), .D (n_1762), .Q
       (n_6447));
  DFRQX1 \integer_file_reg[27][10] (.C (rc_gclk_199975), .D (n_20), .Q
       (n_6788));
  DFRQX1 \integer_file_reg[27][11] (.C (rc_gclk_199975), .D (n_112), .Q
       (n_6819));
  DFRQX1 \integer_file_reg[27][12] (.C (rc_gclk_199975), .D (n_1761),
       .Q (n_6850));
  DFRQX1 \integer_file_reg[27][13] (.C (rc_gclk_199975), .D (n_84), .Q
       (n_6912));
  DFRQX1 \integer_file_reg[27][14] (.C (rc_gclk_199975), .D (n_104), .Q
       (n_6943));
  DFRQX1 \integer_file_reg[27][15] (.C (rc_gclk_199975), .D (n_19), .Q
       (n_6974));
  DFRQX1 \integer_file_reg[27][16] (.C (rc_gclk_199975), .D (n_103), .Q
       (n_7005));
  DFRQX1 \integer_file_reg[27][17] (.C (rc_gclk_199975), .D (n_1760),
       .Q (n_7036));
  DFRQX1 \integer_file_reg[27][18] (.C (rc_gclk_199975), .D (n_22), .Q
       (n_7067));
  DFRQX1 \integer_file_reg[27][19] (.C (rc_gclk_199975), .D (n_1759),
       .Q (n_7098));
  DFRQX1 \integer_file_reg[27][1] (.C (rc_gclk_199975), .D (n_30), .Q
       (n_6478));
  DFRQX1 \integer_file_reg[27][20] (.C (rc_gclk_199975), .D (n_1758),
       .Q (n_7129));
  DFRQX1 \integer_file_reg[27][21] (.C (rc_gclk_199975), .D (n_1757),
       .Q (n_7160));
  DFRQX1 \integer_file_reg[27][22] (.C (rc_gclk_199975), .D (n_1756),
       .Q (n_7191));
  DFRQX1 \integer_file_reg[27][23] (.C (rc_gclk_199975), .D (n_1755),
       .Q (n_6261));
  DFRQX1 \integer_file_reg[27][24] (.C (rc_gclk_199975), .D (n_1754),
       .Q (n_6292));
  DFRQX1 \integer_file_reg[27][25] (.C (rc_gclk_199975), .D (n_1753),
       .Q (n_6323));
  DFRQX1 \integer_file_reg[27][26] (.C (rc_gclk_199975), .D (n_12), .Q
       (n_6354));
  DFRQX1 \integer_file_reg[27][27] (.C (rc_gclk_199975), .D (n_1752),
       .Q (n_6385));
  DFRQX1 \integer_file_reg[27][28] (.C (rc_gclk_199975), .D (n_1751),
       .Q (n_6416));
  DFRQX1 \integer_file_reg[27][29] (.C (rc_gclk_199975), .D (n_1750),
       .Q (n_6540));
  DFRQX1 \integer_file_reg[27][2] (.C (rc_gclk_199975), .D (n_39), .Q
       (n_6509));
  DFRQX1 \integer_file_reg[27][30] (.C (rc_gclk_199975), .D (n_1749),
       .Q (n_6881));
  DFRQX1 \integer_file_reg[27][31] (.C (rc_gclk_199975), .D (n_1748),
       .Q (n_7222));
  DFRQX1 \integer_file_reg[27][3] (.C (rc_gclk_199975), .D (n_25), .Q
       (n_6571));
  DFRQX1 \integer_file_reg[27][4] (.C (rc_gclk_199975), .D (n_51), .Q
       (n_6602));
  DFRQX1 \integer_file_reg[27][5] (.C (rc_gclk_199975), .D (n_49), .Q
       (n_6633));
  DFRQX1 \integer_file_reg[27][6] (.C (rc_gclk_199975), .D (n_46), .Q
       (n_6664));
  DFRQX1 \integer_file_reg[27][7] (.C (rc_gclk_199975), .D (n_81), .Q
       (n_6695));
  DFRQX1 \integer_file_reg[27][8] (.C (rc_gclk_199975), .D (n_101), .Q
       (n_6726));
  DFRQX1 \integer_file_reg[27][9] (.C (rc_gclk_199975), .D (n_100), .Q
       (n_6757));
  DFRQX1 \integer_file_reg[28][0] (.C (rc_gclk_199981), .D (n_1747), .Q
       (n_6446));
  DFRQX1 \integer_file_reg[28][10] (.C (rc_gclk_199981), .D (n_20), .Q
       (n_6787));
  DFRQX1 \integer_file_reg[28][11] (.C (rc_gclk_199981), .D (n_113), .Q
       (n_6818));
  DFRQX1 \integer_file_reg[28][12] (.C (rc_gclk_199981), .D (n_79), .Q
       (n_6849));
  DFRQX1 \integer_file_reg[28][13] (.C (rc_gclk_199981), .D (n_76), .Q
       (n_6911));
  DFRQX1 \integer_file_reg[28][14] (.C (rc_gclk_199981), .D (n_104), .Q
       (n_6942));
  DFRQX1 \integer_file_reg[28][15] (.C (rc_gclk_199981), .D (n_17), .Q
       (n_6973));
  DFRQX1 \integer_file_reg[28][16] (.C (rc_gclk_199981), .D (n_103), .Q
       (n_7004));
  DFRQX1 \integer_file_reg[28][17] (.C (rc_gclk_199981), .D (n_1746),
       .Q (n_7035));
  DFRQX1 \integer_file_reg[28][18] (.C (rc_gclk_199981), .D (n_63), .Q
       (n_7066));
  DFRQX1 \integer_file_reg[28][19] (.C (rc_gclk_199981), .D (n_1745),
       .Q (n_7097));
  DFRQX1 \integer_file_reg[28][1] (.C (rc_gclk_199981), .D (n_30), .Q
       (n_6477));
  DFRQX1 \integer_file_reg[28][20] (.C (rc_gclk_199981), .D (n_1744),
       .Q (n_7128));
  DFRQX1 \integer_file_reg[28][21] (.C (rc_gclk_199981), .D (n_1743),
       .Q (n_7159));
  DFRQX1 \integer_file_reg[28][22] (.C (rc_gclk_199981), .D (n_1742),
       .Q (n_7190));
  DFRQX1 \integer_file_reg[28][23] (.C (rc_gclk_199981), .D (n_1741),
       .Q (n_6260));
  DFRQX1 \integer_file_reg[28][24] (.C (rc_gclk_199981), .D (n_42), .Q
       (n_6291));
  DFRQX1 \integer_file_reg[28][25] (.C (rc_gclk_199981), .D (n_1740),
       .Q (n_6322));
  DFRQX1 \integer_file_reg[28][26] (.C (rc_gclk_199981), .D (n_12), .Q
       (n_6353));
  DFRQX1 \integer_file_reg[28][27] (.C (rc_gclk_199981), .D (n_1739),
       .Q (n_6384));
  DFRQX1 \integer_file_reg[28][28] (.C (rc_gclk_199981), .D (n_1738),
       .Q (n_6415));
  DFRQX1 \integer_file_reg[28][29] (.C (rc_gclk_199981), .D (n_1737),
       .Q (n_6539));
  DFRQX1 \integer_file_reg[28][2] (.C (rc_gclk_199981), .D (n_21), .Q
       (n_6508));
  DFRQX1 \integer_file_reg[28][30] (.C (rc_gclk_199981), .D (n_1736),
       .Q (n_6880));
  DFRQX1 \integer_file_reg[28][31] (.C (rc_gclk_199981), .D (n_1735),
       .Q (n_7221));
  DFRQX1 \integer_file_reg[28][3] (.C (rc_gclk_199981), .D (n_38), .Q
       (n_6570));
  DFRQX1 \integer_file_reg[28][4] (.C (rc_gclk_199981), .D (n_51), .Q
       (n_6601));
  DFRQX1 \integer_file_reg[28][5] (.C (rc_gclk_199981), .D (n_49), .Q
       (n_6632));
  DFRQX1 \integer_file_reg[28][6] (.C (rc_gclk_199981), .D (n_46), .Q
       (n_6663));
  DFRQX1 \integer_file_reg[28][7] (.C (rc_gclk_199981), .D (n_82), .Q
       (n_6694));
  DFRQX1 \integer_file_reg[28][8] (.C (rc_gclk_199981), .D (n_101), .Q
       (n_6725));
  DFRQX1 \integer_file_reg[28][9] (.C (rc_gclk_199981), .D (n_89), .Q
       (n_6756));
  DFRQX1 \integer_file_reg[29][0] (.C (rc_gclk_199984), .D (n_1734), .Q
       (n_6445));
  DFRQX1 \integer_file_reg[29][10] (.C (rc_gclk_199984), .D (n_69), .Q
       (n_6786));
  DFRQX1 \integer_file_reg[29][11] (.C (rc_gclk_199984), .D (n_110), .Q
       (n_6817));
  DFRQX1 \integer_file_reg[29][12] (.C (rc_gclk_199984), .D (n_79), .Q
       (n_6848));
  DFRQX1 \integer_file_reg[29][13] (.C (rc_gclk_199984), .D (n_76), .Q
       (n_6910));
  DFRQX1 \integer_file_reg[29][14] (.C (rc_gclk_199984), .D (n_104), .Q
       (n_6941));
  DFRQX1 \integer_file_reg[29][15] (.C (rc_gclk_199984), .D (n_17), .Q
       (n_6972));
  DFRQX1 \integer_file_reg[29][16] (.C (rc_gclk_199984), .D (n_75), .Q
       (n_7003));
  DFRQX1 \integer_file_reg[29][17] (.C (rc_gclk_199984), .D (n_97), .Q
       (n_7034));
  DFRQX1 \integer_file_reg[29][18] (.C (rc_gclk_199984), .D (n_63), .Q
       (n_7065));
  DFRQX1 \integer_file_reg[29][19] (.C (rc_gclk_199984), .D (n_1733),
       .Q (n_7096));
  DFRQX1 \integer_file_reg[29][1] (.C (rc_gclk_199984), .D (n_26), .Q
       (n_6476));
  DFRQX1 \integer_file_reg[29][20] (.C (rc_gclk_199984), .D (n_1732),
       .Q (n_7127));
  DFRQX1 \integer_file_reg[29][21] (.C (rc_gclk_199984), .D (n_1731),
       .Q (n_7158));
  DFRQX1 \integer_file_reg[29][22] (.C (rc_gclk_199984), .D (n_1730),
       .Q (n_7189));
  DFRQX1 \integer_file_reg[29][23] (.C (rc_gclk_199984), .D (n_1729),
       .Q (n_6259));
  DFRQX1 \integer_file_reg[29][24] (.C (rc_gclk_199984), .D (n_43), .Q
       (n_6290));
  DFRQX1 \integer_file_reg[29][25] (.C (rc_gclk_199984), .D (n_1728),
       .Q (n_6321));
  DFRQX1 \integer_file_reg[29][26] (.C (rc_gclk_199984), .D (n_13), .Q
       (n_6352));
  DFRQX1 \integer_file_reg[29][27] (.C (rc_gclk_199984), .D (n_1727),
       .Q (n_6383));
  DFRQX1 \integer_file_reg[29][28] (.C (rc_gclk_199984), .D (n_1726),
       .Q (n_6414));
  DFRQX1 \integer_file_reg[29][29] (.C (rc_gclk_199984), .D (n_1725),
       .Q (n_6538));
  DFRQX1 \integer_file_reg[29][2] (.C (rc_gclk_199984), .D (n_21), .Q
       (n_6507));
  DFRQX1 \integer_file_reg[29][30] (.C (rc_gclk_199984), .D (n_1724),
       .Q (n_6879));
  DFRQX1 \integer_file_reg[29][31] (.C (rc_gclk_199984), .D (n_1723),
       .Q (n_7220));
  DFRQX1 \integer_file_reg[29][3] (.C (rc_gclk_199984), .D (n_25), .Q
       (n_6569));
  DFRQX1 \integer_file_reg[29][4] (.C (rc_gclk_199984), .D (n_33), .Q
       (n_6600));
  DFRQX1 \integer_file_reg[29][5] (.C (rc_gclk_199984), .D (n_31), .Q
       (n_6631));
  DFRQX1 \integer_file_reg[29][6] (.C (rc_gclk_199984), .D (n_46), .Q
       (n_6662));
  DFRQX1 \integer_file_reg[29][7] (.C (rc_gclk_199984), .D (n_82), .Q
       (n_6693));
  DFRQX1 \integer_file_reg[29][8] (.C (rc_gclk_199984), .D (n_72), .Q
       (n_6724));
  DFRQX1 \integer_file_reg[29][9] (.C (rc_gclk_199984), .D (n_89), .Q
       (n_6755));
  DFRQX1 \integer_file_reg[2][0] (.C (rc_gclk_199891), .D (n_1722), .Q
       (n_6472));
  DFRQX1 \integer_file_reg[2][10] (.C (rc_gclk_199891), .D (n_69), .Q
       (n_6813));
  DFRQX1 \integer_file_reg[2][11] (.C (rc_gclk_199891), .D (n_111), .Q
       (n_6844));
  DFRQX1 \integer_file_reg[2][12] (.C (rc_gclk_199891), .D (n_1721), .Q
       (n_6875));
  DFRQX1 \integer_file_reg[2][13] (.C (rc_gclk_199891), .D (n_76), .Q
       (n_6937));
  DFRQX1 \integer_file_reg[2][14] (.C (rc_gclk_199891), .D (n_104), .Q
       (n_6968));
  DFRQX1 \integer_file_reg[2][15] (.C (rc_gclk_199891), .D (n_18), .Q
       (n_6999));
  DFRQX1 \integer_file_reg[2][16] (.C (rc_gclk_199891), .D (n_75), .Q
       (n_7030));
  DFRQX1 \integer_file_reg[2][17] (.C (rc_gclk_199891), .D (n_1720), .Q
       (n_7061));
  DFRQX1 \integer_file_reg[2][18] (.C (rc_gclk_199891), .D (n_64), .Q
       (n_7092));
  DFRQX1 \integer_file_reg[2][19] (.C (rc_gclk_199891), .D (n_1719), .Q
       (n_7123));
  DFRQX1 \integer_file_reg[2][1] (.C (rc_gclk_199891), .D (n_26), .Q
       (n_6503));
  DFRQX1 \integer_file_reg[2][20] (.C (rc_gclk_199891), .D (n_1718), .Q
       (n_7154));
  DFRQX1 \integer_file_reg[2][21] (.C (rc_gclk_199891), .D (n_1717), .Q
       (n_7185));
  DFRQX1 \integer_file_reg[2][22] (.C (rc_gclk_199891), .D (n_1716), .Q
       (n_7216));
  DFRQX1 \integer_file_reg[2][23] (.C (rc_gclk_199891), .D (n_1715), .Q
       (n_6286));
  DFRQX1 \integer_file_reg[2][24] (.C (rc_gclk_199891), .D (n_1714), .Q
       (n_6317));
  DFRQX1 \integer_file_reg[2][25] (.C (rc_gclk_199891), .D (n_1713), .Q
       (n_6348));
  DFRQX1 \integer_file_reg[2][26] (.C (rc_gclk_199891), .D (n_13), .Q
       (n_6379));
  DFRQX1 \integer_file_reg[2][27] (.C (rc_gclk_199891), .D (n_1712), .Q
       (n_6410));
  DFRQX1 \integer_file_reg[2][28] (.C (rc_gclk_199891), .D (n_1711), .Q
       (n_6441));
  DFRQX1 \integer_file_reg[2][29] (.C (rc_gclk_199891), .D (n_1710), .Q
       (n_6565));
  DFRQX1 \integer_file_reg[2][2] (.C (rc_gclk_199891), .D (n_21), .Q
       (n_6534));
  DFRQX1 \integer_file_reg[2][30] (.C (rc_gclk_199891), .D (n_1709), .Q
       (n_6906));
  DFRQX1 \integer_file_reg[2][31] (.C (rc_gclk_199891), .D (n_1708), .Q
       (n_7247));
  DFRQX1 \integer_file_reg[2][3] (.C (rc_gclk_199891), .D (n_53), .Q
       (n_6596));
  DFRQX1 \integer_file_reg[2][4] (.C (rc_gclk_199891), .D (n_28), .Q
       (n_6627));
  DFRQX1 \integer_file_reg[2][5] (.C (rc_gclk_199891), .D (n_32), .Q
       (n_6658));
  DFRQX1 \integer_file_reg[2][6] (.C (rc_gclk_199891), .D (n_27), .Q
       (n_6689));
  DFRQX1 \integer_file_reg[2][7] (.C (rc_gclk_199891), .D (n_82), .Q
       (n_6720));
  DFRQX1 \integer_file_reg[2][8] (.C (rc_gclk_199891), .D (n_72), .Q
       (n_6751));
  DFRQX1 \integer_file_reg[2][9] (.C (rc_gclk_199891), .D (n_89), .Q
       (n_6782));
  DFRQX1 \integer_file_reg[30][0] (.C (rc_gclk_199894), .D (n_1707), .Q
       (n_6444));
  DFRQX1 \integer_file_reg[30][10] (.C (rc_gclk_199894), .D (n_20), .Q
       (n_6785));
  DFRQX1 \integer_file_reg[30][11] (.C (rc_gclk_199894), .D (n_110), .Q
       (n_6816));
  DFRQX1 \integer_file_reg[30][12] (.C (rc_gclk_199894), .D (n_1706),
       .Q (n_6847));
  DFRQX1 \integer_file_reg[30][13] (.C (rc_gclk_199894), .D (n_76), .Q
       (n_6909));
  DFRQX1 \integer_file_reg[30][14] (.C (rc_gclk_199894), .D (n_71), .Q
       (n_6940));
  DFRQX1 \integer_file_reg[30][15] (.C (rc_gclk_199894), .D (n_18), .Q
       (n_6971));
  DFRQX1 \integer_file_reg[30][16] (.C (rc_gclk_199894), .D (n_75), .Q
       (n_7002));
  DFRQX1 \integer_file_reg[30][17] (.C (rc_gclk_199894), .D (n_1705),
       .Q (n_7033));
  DFRQX1 \integer_file_reg[30][18] (.C (rc_gclk_199894), .D (n_64), .Q
       (n_7064));
  DFRQX1 \integer_file_reg[30][19] (.C (rc_gclk_199894), .D (n_1704),
       .Q (n_7095));
  DFRQX1 \integer_file_reg[30][1] (.C (rc_gclk_199894), .D (n_24), .Q
       (n_6475));
  DFRQX1 \integer_file_reg[30][20] (.C (rc_gclk_199894), .D (n_1703),
       .Q (n_7126));
  DFRQX1 \integer_file_reg[30][21] (.C (rc_gclk_199894), .D (n_1702),
       .Q (n_7157));
  DFRQX1 \integer_file_reg[30][22] (.C (rc_gclk_199894), .D (n_1701),
       .Q (n_7188));
  DFRQX1 \integer_file_reg[30][23] (.C (rc_gclk_199894), .D (n_1700),
       .Q (n_6258));
  DFRQX1 \integer_file_reg[30][24] (.C (rc_gclk_199894), .D (n_43), .Q
       (n_6289));
  DFRQX1 \integer_file_reg[30][25] (.C (rc_gclk_199894), .D (n_1699),
       .Q (n_6320));
  DFRQX1 \integer_file_reg[30][26] (.C (rc_gclk_199894), .D (n_14), .Q
       (n_6351));
  DFRQX1 \integer_file_reg[30][27] (.C (rc_gclk_199894), .D (n_1698),
       .Q (n_6382));
  DFRQX1 \integer_file_reg[30][28] (.C (rc_gclk_199894), .D (n_1697),
       .Q (n_6413));
  DFRQX1 \integer_file_reg[30][29] (.C (rc_gclk_199894), .D (n_1696),
       .Q (n_6537));
  DFRQX1 \integer_file_reg[30][2] (.C (rc_gclk_199894), .D (n_21), .Q
       (n_6506));
  DFRQX1 \integer_file_reg[30][30] (.C (rc_gclk_199894), .D (n_1695),
       .Q (n_6878));
  DFRQX1 \integer_file_reg[30][31] (.C (rc_gclk_199894), .D (n_1694),
       .Q (n_7219));
  DFRQX1 \integer_file_reg[30][3] (.C (rc_gclk_199894), .D (n_53), .Q
       (n_6568));
  DFRQX1 \integer_file_reg[30][4] (.C (rc_gclk_199894), .D (n_28), .Q
       (n_6599));
  DFRQX1 \integer_file_reg[30][5] (.C (rc_gclk_199894), .D (n_23), .Q
       (n_6630));
  DFRQX1 \integer_file_reg[30][6] (.C (rc_gclk_199894), .D (n_27), .Q
       (n_6661));
  DFRQX1 \integer_file_reg[30][7] (.C (rc_gclk_199894), .D (n_81), .Q
       (n_6692));
  DFRQX1 \integer_file_reg[30][8] (.C (rc_gclk_199894), .D (n_72), .Q
       (n_6723));
  DFRQX1 \integer_file_reg[30][9] (.C (rc_gclk_199894), .D (n_89), .Q
       (n_6754));
  DFRQX1 \integer_file_reg[31][0] (.C (rc_gclk_199900), .D (n_1693), .Q
       (n_6443));
  DFRQX1 \integer_file_reg[31][10] (.C (rc_gclk_199900), .D (n_20), .Q
       (n_6784));
  DFRQX1 \integer_file_reg[31][11] (.C (rc_gclk_199900), .D (n_112), .Q
       (n_6815));
  DFRQX1 \integer_file_reg[31][12] (.C (rc_gclk_199900), .D (n_1692),
       .Q (n_6846));
  DFRQX1 \integer_file_reg[31][13] (.C (rc_gclk_199900), .D (n_76), .Q
       (n_6908));
  DFRQX1 \integer_file_reg[31][14] (.C (rc_gclk_199900), .D (n_71), .Q
       (n_6939));
  DFRQX1 \integer_file_reg[31][15] (.C (rc_gclk_199900), .D (n_18), .Q
       (n_6970));
  DFRQX1 \integer_file_reg[31][16] (.C (rc_gclk_199900), .D (n_75), .Q
       (n_7001));
  DFRQX1 \integer_file_reg[31][17] (.C (rc_gclk_199900), .D (n_91), .Q
       (n_7032));
  DFRQX1 \integer_file_reg[31][18] (.C (rc_gclk_199900), .D (n_65), .Q
       (n_7063));
  DFRQX1 \integer_file_reg[31][19] (.C (rc_gclk_199900), .D (n_1691),
       .Q (n_7094));
  DFRQX1 \integer_file_reg[31][1] (.C (rc_gclk_199900), .D (n_24), .Q
       (n_6474));
  DFRQX1 \integer_file_reg[31][20] (.C (rc_gclk_199900), .D (n_1690),
       .Q (n_7125));
  DFRQX1 \integer_file_reg[31][21] (.C (rc_gclk_199900), .D (n_1689),
       .Q (n_7156));
  DFRQX1 \integer_file_reg[31][22] (.C (rc_gclk_199900), .D (n_1688),
       .Q (n_7187));
  DFRQX1 \integer_file_reg[31][23] (.C (rc_gclk_199900), .D (n_1687),
       .Q (n_6257));
  DFRQX1 \integer_file_reg[31][24] (.C (rc_gclk_199900), .D (n_44), .Q
       (n_6288));
  DFRQX1 \integer_file_reg[31][25] (.C (rc_gclk_199900), .D (n_1686),
       .Q (n_6319));
  DFRQX1 \integer_file_reg[31][26] (.C (rc_gclk_199900), .D (n_14), .Q
       (n_6350));
  DFRQX1 \integer_file_reg[31][27] (.C (rc_gclk_199900), .D (n_1685),
       .Q (n_6381));
  DFRQX1 \integer_file_reg[31][28] (.C (rc_gclk_199900), .D (n_1684),
       .Q (n_6412));
  DFRQX1 \integer_file_reg[31][29] (.C (rc_gclk_199900), .D (n_1683),
       .Q (n_6536));
  DFRQX1 \integer_file_reg[31][2] (.C (rc_gclk_199900), .D (n_54), .Q
       (n_6505));
  DFRQX1 \integer_file_reg[31][30] (.C (rc_gclk_199900), .D (n_1682),
       .Q (n_6877));
  DFRQX1 \integer_file_reg[31][31] (.C (rc_gclk_199900), .D (n_1681),
       .Q (n_7218));
  DFRQX1 \integer_file_reg[31][3] (.C (rc_gclk_199900), .D (n_25), .Q
       (n_6567));
  DFRQX1 \integer_file_reg[31][4] (.C (rc_gclk_199900), .D (n_29), .Q
       (n_6598));
  DFRQX1 \integer_file_reg[31][5] (.C (rc_gclk_199900), .D (n_23), .Q
       (n_6629));
  DFRQX1 \integer_file_reg[31][6] (.C (rc_gclk_199900), .D (n_46), .Q
       (n_6660));
  DFRQX1 \integer_file_reg[31][7] (.C (rc_gclk_199900), .D (n_81), .Q
       (n_6691));
  DFRQX1 \integer_file_reg[31][8] (.C (rc_gclk_199900), .D (n_72), .Q
       (n_6722));
  DFRQX1 \integer_file_reg[31][9] (.C (rc_gclk_199900), .D (n_78), .Q
       (n_6753));
  DFRQX1 \integer_file_reg[3][0] (.C (rc_gclk_199903), .D (n_1680), .Q
       (n_6471));
  DFRQX1 \integer_file_reg[3][10] (.C (rc_gclk_199903), .D (n_69), .Q
       (n_6812));
  DFRQX1 \integer_file_reg[3][11] (.C (rc_gclk_199903), .D (n_113), .Q
       (n_6843));
  DFRQX1 \integer_file_reg[3][12] (.C (rc_gclk_199903), .D (n_1679), .Q
       (n_6874));
  DFRQX1 \integer_file_reg[3][13] (.C (rc_gclk_199903), .D (n_76), .Q
       (n_6936));
  DFRQX1 \integer_file_reg[3][14] (.C (rc_gclk_199903), .D (n_71), .Q
       (n_6967));
  DFRQX1 \integer_file_reg[3][15] (.C (rc_gclk_199903), .D (n_18), .Q
       (n_6998));
  DFRQX1 \integer_file_reg[3][16] (.C (rc_gclk_199903), .D (n_98), .Q
       (n_7029));
  DFRQX1 \integer_file_reg[3][17] (.C (rc_gclk_199903), .D (n_91), .Q
       (n_7060));
  DFRQX1 \integer_file_reg[3][18] (.C (rc_gclk_199903), .D (n_65), .Q
       (n_7091));
  DFRQX1 \integer_file_reg[3][19] (.C (rc_gclk_199903), .D (n_1678), .Q
       (n_7122));
  DFRQX1 \integer_file_reg[3][1] (.C (rc_gclk_199903), .D (n_26), .Q
       (n_6502));
  DFRQX1 \integer_file_reg[3][20] (.C (rc_gclk_199903), .D (n_1677), .Q
       (n_7153));
  DFRQX1 \integer_file_reg[3][21] (.C (rc_gclk_199903), .D (n_1676), .Q
       (n_7184));
  DFRQX1 \integer_file_reg[3][22] (.C (rc_gclk_199903), .D (n_1675), .Q
       (n_7215));
  DFRQX1 \integer_file_reg[3][23] (.C (rc_gclk_199903), .D (n_1674), .Q
       (n_6285));
  DFRQX1 \integer_file_reg[3][24] (.C (rc_gclk_199903), .D (n_1673), .Q
       (n_6316));
  DFRQX1 \integer_file_reg[3][25] (.C (rc_gclk_199903), .D (n_1672), .Q
       (n_6347));
  DFRQX1 \integer_file_reg[3][26] (.C (rc_gclk_199903), .D (n_4), .Q
       (n_6378));
  DFRQX1 \integer_file_reg[3][27] (.C (rc_gclk_199903), .D (n_1671), .Q
       (n_6409));
  DFRQX1 \integer_file_reg[3][28] (.C (rc_gclk_199903), .D (n_1670), .Q
       (n_6440));
  DFRQX1 \integer_file_reg[3][29] (.C (rc_gclk_199903), .D (n_1669), .Q
       (n_6564));
  DFRQX1 \integer_file_reg[3][2] (.C (rc_gclk_199903), .D (n_54), .Q
       (n_6533));
  DFRQX1 \integer_file_reg[3][30] (.C (rc_gclk_199903), .D (n_1668), .Q
       (n_6905));
  DFRQX1 \integer_file_reg[3][31] (.C (rc_gclk_199903), .D (n_1667), .Q
       (n_7246));
  DFRQX1 \integer_file_reg[3][3] (.C (rc_gclk_199903), .D (n_38), .Q
       (n_6595));
  DFRQX1 \integer_file_reg[3][4] (.C (rc_gclk_199903), .D (n_29), .Q
       (n_6626));
  DFRQX1 \integer_file_reg[3][5] (.C (rc_gclk_199903), .D (n_31), .Q
       (n_6657));
  DFRQX1 \integer_file_reg[3][6] (.C (rc_gclk_199903), .D (n_46), .Q
       (n_6688));
  DFRQX1 \integer_file_reg[3][7] (.C (rc_gclk_199903), .D (n_82), .Q
       (n_6719));
  DFRQX1 \integer_file_reg[3][8] (.C (rc_gclk_199903), .D (n_101), .Q
       (n_6750));
  DFRQX1 \integer_file_reg[3][9] (.C (rc_gclk_199903), .D (n_100), .Q
       (n_6781));
  DFRQX1 \integer_file_reg[4][0] (.C (rc_gclk_199909), .D (n_1666), .Q
       (n_6470));
  DFRQX1 \integer_file_reg[4][10] (.C (rc_gclk_199909), .D (n_69), .Q
       (n_6811));
  DFRQX1 \integer_file_reg[4][11] (.C (rc_gclk_199909), .D (n_111), .Q
       (n_6842));
  DFRQX1 \integer_file_reg[4][12] (.C (rc_gclk_199909), .D (n_1665), .Q
       (n_6873));
  DFRQX1 \integer_file_reg[4][13] (.C (rc_gclk_199909), .D (n_88), .Q
       (n_6935));
  DFRQX1 \integer_file_reg[4][14] (.C (rc_gclk_199909), .D (n_71), .Q
       (n_6966));
  DFRQX1 \integer_file_reg[4][15] (.C (rc_gclk_199909), .D (n_17), .Q
       (n_6997));
  DFRQX1 \integer_file_reg[4][16] (.C (rc_gclk_199909), .D (n_98), .Q
       (n_7028));
  DFRQX1 \integer_file_reg[4][17] (.C (rc_gclk_199909), .D (n_91), .Q
       (n_7059));
  DFRQX1 \integer_file_reg[4][18] (.C (rc_gclk_199909), .D (n_66), .Q
       (n_7090));
  DFRQX1 \integer_file_reg[4][19] (.C (rc_gclk_199909), .D (n_1664), .Q
       (n_7121));
  DFRQX1 \integer_file_reg[4][1] (.C (rc_gclk_199909), .D (n_26), .Q
       (n_6501));
  DFRQX1 \integer_file_reg[4][20] (.C (rc_gclk_199909), .D (n_1663), .Q
       (n_7152));
  DFRQX1 \integer_file_reg[4][21] (.C (rc_gclk_199909), .D (n_1662), .Q
       (n_7183));
  DFRQX1 \integer_file_reg[4][22] (.C (rc_gclk_199909), .D (n_1661), .Q
       (n_7214));
  DFRQX1 \integer_file_reg[4][23] (.C (rc_gclk_199909), .D (n_1660), .Q
       (n_6284));
  DFRQX1 \integer_file_reg[4][24] (.C (rc_gclk_199909), .D (n_1659), .Q
       (n_6315));
  DFRQX1 \integer_file_reg[4][25] (.C (rc_gclk_199909), .D (n_1658), .Q
       (n_6346));
  DFRQX1 \integer_file_reg[4][26] (.C (rc_gclk_199909), .D (n_5), .Q
       (n_6377));
  DFRQX1 \integer_file_reg[4][27] (.C (rc_gclk_199909), .D (n_1657), .Q
       (n_6408));
  DFRQX1 \integer_file_reg[4][28] (.C (rc_gclk_199909), .D (n_1656), .Q
       (n_6439));
  DFRQX1 \integer_file_reg[4][29] (.C (rc_gclk_199909), .D (n_1655), .Q
       (n_6563));
  DFRQX1 \integer_file_reg[4][2] (.C (rc_gclk_199909), .D (n_54), .Q
       (n_6532));
  DFRQX1 \integer_file_reg[4][30] (.C (rc_gclk_199909), .D (n_1654), .Q
       (n_6904));
  DFRQX1 \integer_file_reg[4][31] (.C (rc_gclk_199909), .D (n_1653), .Q
       (n_7245));
  DFRQX1 \integer_file_reg[4][3] (.C (rc_gclk_199909), .D (n_38), .Q
       (n_6594));
  DFRQX1 \integer_file_reg[4][4] (.C (rc_gclk_199909), .D (n_28), .Q
       (n_6625));
  DFRQX1 \integer_file_reg[4][5] (.C (rc_gclk_199909), .D (n_32), .Q
       (n_6656));
  DFRQX1 \integer_file_reg[4][6] (.C (rc_gclk_199909), .D (n_37), .Q
       (n_6687));
  DFRQX1 \integer_file_reg[4][7] (.C (rc_gclk_199909), .D (n_81), .Q
       (n_6718));
  DFRQX1 \integer_file_reg[4][8] (.C (rc_gclk_199909), .D (n_101), .Q
       (n_6749));
  DFRQX1 \integer_file_reg[4][9] (.C (rc_gclk_199909), .D (n_89), .Q
       (n_6780));
  DFRQX1 \integer_file_reg[5][0] (.C (rc_gclk_199912), .D (n_1652), .Q
       (n_6469));
  DFRQX1 \integer_file_reg[5][10] (.C (rc_gclk_199912), .D (n_20), .Q
       (n_6810));
  DFRQX1 \integer_file_reg[5][11] (.C (rc_gclk_199912), .D (n_110), .Q
       (n_6841));
  DFRQX1 \integer_file_reg[5][12] (.C (rc_gclk_199912), .D (n_1651), .Q
       (n_6872));
  DFRQX1 \integer_file_reg[5][13] (.C (rc_gclk_199912), .D (n_76), .Q
       (n_6934));
  DFRQX1 \integer_file_reg[5][14] (.C (rc_gclk_199912), .D (n_73), .Q
       (n_6965));
  DFRQX1 \integer_file_reg[5][15] (.C (rc_gclk_199912), .D (n_17), .Q
       (n_6996));
  DFRQX1 \integer_file_reg[5][16] (.C (rc_gclk_199912), .D (n_75), .Q
       (n_7027));
  DFRQX1 \integer_file_reg[5][17] (.C (rc_gclk_199912), .D (n_91), .Q
       (n_7058));
  DFRQX1 \integer_file_reg[5][18] (.C (rc_gclk_199912), .D (n_66), .Q
       (n_7089));
  DFRQX1 \integer_file_reg[5][19] (.C (rc_gclk_199912), .D (n_1650), .Q
       (n_7120));
  DFRQX1 \integer_file_reg[5][1] (.C (rc_gclk_199912), .D (n_24), .Q
       (n_6500));
  DFRQX1 \integer_file_reg[5][20] (.C (rc_gclk_199912), .D (n_1649), .Q
       (n_7151));
  DFRQX1 \integer_file_reg[5][21] (.C (rc_gclk_199912), .D (n_1648), .Q
       (n_7182));
  DFRQX1 \integer_file_reg[5][22] (.C (rc_gclk_199912), .D (n_1647), .Q
       (n_7213));
  DFRQX1 \integer_file_reg[5][23] (.C (rc_gclk_199912), .D (n_1646), .Q
       (n_6283));
  DFRQX1 \integer_file_reg[5][24] (.C (rc_gclk_199912), .D (n_1645), .Q
       (n_6314));
  DFRQX1 \integer_file_reg[5][25] (.C (rc_gclk_199912), .D (n_1644), .Q
       (n_6345));
  DFRQX1 \integer_file_reg[5][26] (.C (rc_gclk_199912), .D (n_15), .Q
       (n_6376));
  DFRQX1 \integer_file_reg[5][27] (.C (rc_gclk_199912), .D (n_1643), .Q
       (n_6407));
  DFRQX1 \integer_file_reg[5][28] (.C (rc_gclk_199912), .D (n_1642), .Q
       (n_6438));
  DFRQX1 \integer_file_reg[5][29] (.C (rc_gclk_199912), .D (n_1641), .Q
       (n_6562));
  DFRQX1 \integer_file_reg[5][2] (.C (rc_gclk_199912), .D (n_54), .Q
       (n_6531));
  DFRQX1 \integer_file_reg[5][30] (.C (rc_gclk_199912), .D (n_1640), .Q
       (n_6903));
  DFRQX1 \integer_file_reg[5][31] (.C (rc_gclk_199912), .D (n_1639), .Q
       (n_7244));
  DFRQX1 \integer_file_reg[5][3] (.C (rc_gclk_199912), .D (n_38), .Q
       (n_6593));
  DFRQX1 \integer_file_reg[5][4] (.C (rc_gclk_199912), .D (n_34), .Q
       (n_6624));
  DFRQX1 \integer_file_reg[5][5] (.C (rc_gclk_199912), .D (n_23), .Q
       (n_6655));
  DFRQX1 \integer_file_reg[5][6] (.C (rc_gclk_199912), .D (n_37), .Q
       (n_6686));
  DFRQX1 \integer_file_reg[5][7] (.C (rc_gclk_199912), .D (n_82), .Q
       (n_6717));
  DFRQX1 \integer_file_reg[5][8] (.C (rc_gclk_199912), .D (n_80), .Q
       (n_6748));
  DFRQX1 \integer_file_reg[5][9] (.C (rc_gclk_199912), .D (n_99), .Q
       (n_6779));
  DFRQX1 \integer_file_reg[6][0] (.C (rc_gclk_199918), .D (n_1638), .Q
       (n_6468));
  DFRQX1 \integer_file_reg[6][10] (.C (rc_gclk_199918), .D (n_20), .Q
       (n_6809));
  DFRQX1 \integer_file_reg[6][11] (.C (rc_gclk_199918), .D (n_113), .Q
       (n_6840));
  DFRQX1 \integer_file_reg[6][12] (.C (rc_gclk_199918), .D (n_79), .Q
       (n_6871));
  DFRQX1 \integer_file_reg[6][13] (.C (rc_gclk_199918), .D (n_106), .Q
       (n_6933));
  DFRQX1 \integer_file_reg[6][14] (.C (rc_gclk_199918), .D (n_73), .Q
       (n_6964));
  DFRQX1 \integer_file_reg[6][15] (.C (rc_gclk_199918), .D (n_19), .Q
       (n_6995));
  DFRQX1 \integer_file_reg[6][16] (.C (rc_gclk_199918), .D (n_75), .Q
       (n_7026));
  DFRQX1 \integer_file_reg[6][17] (.C (rc_gclk_199918), .D (n_1637), .Q
       (n_7057));
  DFRQX1 \integer_file_reg[6][18] (.C (rc_gclk_199918), .D (n_67), .Q
       (n_7088));
  DFRQX1 \integer_file_reg[6][19] (.C (rc_gclk_199918), .D (n_1636), .Q
       (n_7119));
  DFRQX1 \integer_file_reg[6][1] (.C (rc_gclk_199918), .D (n_24), .Q
       (n_6499));
  DFRQX1 \integer_file_reg[6][20] (.C (rc_gclk_199918), .D (n_1635), .Q
       (n_7150));
  DFRQX1 \integer_file_reg[6][21] (.C (rc_gclk_199918), .D (n_1634), .Q
       (n_7181));
  DFRQX1 \integer_file_reg[6][22] (.C (rc_gclk_199918), .D (n_1633), .Q
       (n_7212));
  DFRQX1 \integer_file_reg[6][23] (.C (rc_gclk_199918), .D (n_1632), .Q
       (n_6282));
  DFRQX1 \integer_file_reg[6][24] (.C (rc_gclk_199918), .D (n_1631), .Q
       (n_6313));
  DFRQX1 \integer_file_reg[6][25] (.C (rc_gclk_199918), .D (n_1630), .Q
       (n_6344));
  DFRQX1 \integer_file_reg[6][26] (.C (rc_gclk_199918), .D (n_15), .Q
       (n_6375));
  DFRQX1 \integer_file_reg[6][27] (.C (rc_gclk_199918), .D (n_1629), .Q
       (n_6406));
  DFRQX1 \integer_file_reg[6][28] (.C (rc_gclk_199918), .D (n_1628), .Q
       (n_6437));
  DFRQX1 \integer_file_reg[6][29] (.C (rc_gclk_199918), .D (n_1627), .Q
       (n_6561));
  DFRQX1 \integer_file_reg[6][2] (.C (rc_gclk_199918), .D (n_39), .Q
       (n_6530));
  DFRQX1 \integer_file_reg[6][30] (.C (rc_gclk_199918), .D (n_1626), .Q
       (n_6902));
  DFRQX1 \integer_file_reg[6][31] (.C (rc_gclk_199918), .D (n_1625), .Q
       (n_7243));
  DFRQX1 \integer_file_reg[6][3] (.C (rc_gclk_199918), .D (n_25), .Q
       (n_6592));
  DFRQX1 \integer_file_reg[6][4] (.C (rc_gclk_199918), .D (n_35), .Q
       (n_6623));
  DFRQX1 \integer_file_reg[6][5] (.C (rc_gclk_199918), .D (n_23), .Q
       (n_6654));
  DFRQX1 \integer_file_reg[6][6] (.C (rc_gclk_199918), .D (n_46), .Q
       (n_6685));
  DFRQX1 \integer_file_reg[6][7] (.C (rc_gclk_199918), .D (n_82), .Q
       (n_6716));
  DFRQX1 \integer_file_reg[6][8] (.C (rc_gclk_199918), .D (n_80), .Q
       (n_6747));
  DFRQX1 \integer_file_reg[6][9] (.C (rc_gclk_199918), .D (n_89), .Q
       (n_6778));
  DFRQX1 \integer_file_reg[7][0] (.C (rc_gclk_199921), .D (n_1624), .Q
       (n_6467));
  DFRQX1 \integer_file_reg[7][10] (.C (rc_gclk_199921), .D (n_69), .Q
       (n_6808));
  DFRQX1 \integer_file_reg[7][11] (.C (rc_gclk_199921), .D (n_110), .Q
       (n_6839));
  DFRQX1 \integer_file_reg[7][12] (.C (rc_gclk_199921), .D (n_77), .Q
       (n_6870));
  DFRQX1 \integer_file_reg[7][13] (.C (rc_gclk_199921), .D (n_109), .Q
       (n_6932));
  DFRQX1 \integer_file_reg[7][14] (.C (rc_gclk_199921), .D (n_73), .Q
       (n_6963));
  DFRQX1 \integer_file_reg[7][15] (.C (rc_gclk_199921), .D (n_19), .Q
       (n_6994));
  DFRQX1 \integer_file_reg[7][16] (.C (rc_gclk_199921), .D (n_98), .Q
       (n_7025));
  DFRQX1 \integer_file_reg[7][17] (.C (rc_gclk_199921), .D (n_91), .Q
       (n_7056));
  DFRQX1 \integer_file_reg[7][18] (.C (rc_gclk_199921), .D (n_67), .Q
       (n_7087));
  DFRQX1 \integer_file_reg[7][19] (.C (rc_gclk_199921), .D (n_1623), .Q
       (n_7118));
  DFRQX1 \integer_file_reg[7][1] (.C (rc_gclk_199921), .D (n_24), .Q
       (n_6498));
  DFRQX1 \integer_file_reg[7][20] (.C (rc_gclk_199921), .D (n_1622), .Q
       (n_7149));
  DFRQX1 \integer_file_reg[7][21] (.C (rc_gclk_199921), .D (n_1621), .Q
       (n_7180));
  DFRQX1 \integer_file_reg[7][22] (.C (rc_gclk_199921), .D (n_1620), .Q
       (n_7211));
  DFRQX1 \integer_file_reg[7][23] (.C (rc_gclk_199921), .D (n_1619), .Q
       (n_6281));
  DFRQX1 \integer_file_reg[7][24] (.C (rc_gclk_199921), .D (n_44), .Q
       (n_6312));
  DFRQX1 \integer_file_reg[7][25] (.C (rc_gclk_199921), .D (n_1618), .Q
       (n_6343));
  DFRQX1 \integer_file_reg[7][26] (.C (rc_gclk_199921), .D (n_5), .Q
       (n_6374));
  DFRQX1 \integer_file_reg[7][27] (.C (rc_gclk_199921), .D (n_1617), .Q
       (n_6405));
  DFRQX1 \integer_file_reg[7][28] (.C (rc_gclk_199921), .D (n_1616), .Q
       (n_6436));
  DFRQX1 \integer_file_reg[7][29] (.C (rc_gclk_199921), .D (n_1615), .Q
       (n_6560));
  DFRQX1 \integer_file_reg[7][2] (.C (rc_gclk_199921), .D (n_39), .Q
       (n_6529));
  DFRQX1 \integer_file_reg[7][30] (.C (rc_gclk_199921), .D (n_1614), .Q
       (n_6901));
  DFRQX1 \integer_file_reg[7][31] (.C (rc_gclk_199921), .D (n_1613), .Q
       (n_7242));
  DFRQX1 \integer_file_reg[7][3] (.C (rc_gclk_199921), .D (n_53), .Q
       (n_6591));
  DFRQX1 \integer_file_reg[7][4] (.C (rc_gclk_199921), .D (n_28), .Q
       (n_6622));
  DFRQX1 \integer_file_reg[7][5] (.C (rc_gclk_199921), .D (n_31), .Q
       (n_6653));
  DFRQX1 \integer_file_reg[7][6] (.C (rc_gclk_199921), .D (n_46), .Q
       (n_6684));
  DFRQX1 \integer_file_reg[7][7] (.C (rc_gclk_199921), .D (n_81), .Q
       (n_6715));
  DFRQX1 \integer_file_reg[7][8] (.C (rc_gclk_199921), .D (n_72), .Q
       (n_6746));
  DFRQX1 \integer_file_reg[7][9] (.C (rc_gclk_199921), .D (n_89), .Q
       (n_6777));
  DFRQX1 \integer_file_reg[8][0] (.C (rc_gclk_199930), .D (n_1612), .Q
       (n_6466));
  DFRQX1 \integer_file_reg[8][10] (.C (rc_gclk_199930), .D (n_70), .Q
       (n_6807));
  DFRQX1 \integer_file_reg[8][11] (.C (rc_gclk_199930), .D (n_110), .Q
       (n_6838));
  DFRQX1 \integer_file_reg[8][12] (.C (rc_gclk_199930), .D (n_77), .Q
       (n_6869));
  DFRQX1 \integer_file_reg[8][13] (.C (rc_gclk_199930), .D (n_107), .Q
       (n_6931));
  DFRQX1 \integer_file_reg[8][14] (.C (rc_gclk_199930), .D (n_71), .Q
       (n_6962));
  DFRQX1 \integer_file_reg[8][15] (.C (rc_gclk_199930), .D (n_17), .Q
       (n_6993));
  DFRQX1 \integer_file_reg[8][16] (.C (rc_gclk_199930), .D (n_75), .Q
       (n_7024));
  DFRQX1 \integer_file_reg[8][17] (.C (rc_gclk_199930), .D (n_91), .Q
       (n_7055));
  DFRQX1 \integer_file_reg[8][18] (.C (rc_gclk_199930), .D (n_68), .Q
       (n_7086));
  DFRQX1 \integer_file_reg[8][19] (.C (rc_gclk_199930), .D (n_1611), .Q
       (n_7117));
  DFRQX1 \integer_file_reg[8][1] (.C (rc_gclk_199930), .D (n_24), .Q
       (n_6497));
  DFRQX1 \integer_file_reg[8][20] (.C (rc_gclk_199930), .D (n_1610), .Q
       (n_7148));
  DFRQX1 \integer_file_reg[8][21] (.C (rc_gclk_199930), .D (n_1609), .Q
       (n_7179));
  DFRQX1 \integer_file_reg[8][22] (.C (rc_gclk_199930), .D (n_1608), .Q
       (n_7210));
  DFRQX1 \integer_file_reg[8][23] (.C (rc_gclk_199930), .D (n_1607), .Q
       (n_6280));
  DFRQX1 \integer_file_reg[8][24] (.C (rc_gclk_199930), .D (n_45), .Q
       (n_6311));
  DFRQX1 \integer_file_reg[8][25] (.C (rc_gclk_199930), .D (n_1606), .Q
       (n_6342));
  DFRQX1 \integer_file_reg[8][26] (.C (rc_gclk_199930), .D (n_16), .Q
       (n_6373));
  DFRQX1 \integer_file_reg[8][27] (.C (rc_gclk_199930), .D (n_1605), .Q
       (n_6404));
  DFRQX1 \integer_file_reg[8][28] (.C (rc_gclk_199930), .D (n_1604), .Q
       (n_6435));
  DFRQX1 \integer_file_reg[8][29] (.C (rc_gclk_199930), .D (n_1603), .Q
       (n_6559));
  DFRQX1 \integer_file_reg[8][2] (.C (rc_gclk_199930), .D (n_54), .Q
       (n_6528));
  DFRQX1 \integer_file_reg[8][30] (.C (rc_gclk_199930), .D (n_1602), .Q
       (n_6900));
  DFRQX1 \integer_file_reg[8][31] (.C (rc_gclk_199930), .D (n_1601), .Q
       (n_7241));
  DFRQX1 \integer_file_reg[8][3] (.C (rc_gclk_199930), .D (n_53), .Q
       (n_6590));
  DFRQX1 \integer_file_reg[8][4] (.C (rc_gclk_199930), .D (n_28), .Q
       (n_6621));
  DFRQX1 \integer_file_reg[8][5] (.C (rc_gclk_199930), .D (n_32), .Q
       (n_6652));
  DFRQX1 \integer_file_reg[8][6] (.C (rc_gclk_199930), .D (n_46), .Q
       (n_6683));
  DFRQX1 \integer_file_reg[8][7] (.C (rc_gclk_199930), .D (n_81), .Q
       (n_6714));
  DFRQX1 \integer_file_reg[8][8] (.C (rc_gclk_199930), .D (n_72), .Q
       (n_6745));
  DFRQX1 \integer_file_reg[8][9] (.C (rc_gclk_199930), .D (n_99), .Q
       (n_6776));
  DFRQX1 \integer_file_reg[9][0] (.C (rc_gclk_199933), .D (n_1600), .Q
       (n_6465));
  DFRQX1 \integer_file_reg[9][10] (.C (rc_gclk_199933), .D (n_70), .Q
       (n_6806));
  DFRQX1 \integer_file_reg[9][11] (.C (rc_gclk_199933), .D (n_112), .Q
       (n_6837));
  DFRQX1 \integer_file_reg[9][12] (.C (rc_gclk_199933), .D (n_77), .Q
       (n_6868));
  DFRQX1 \integer_file_reg[9][13] (.C (rc_gclk_199933), .D (n_83), .Q
       (n_6930));
  DFRQX1 \integer_file_reg[9][14] (.C (rc_gclk_199933), .D (n_71), .Q
       (n_6961));
  DFRQX1 \integer_file_reg[9][15] (.C (rc_gclk_199933), .D (n_17), .Q
       (n_6992));
  DFRQX1 \integer_file_reg[9][16] (.C (rc_gclk_199933), .D (n_98), .Q
       (n_7023));
  DFRQX1 \integer_file_reg[9][17] (.C (rc_gclk_199933), .D (n_1599), .Q
       (n_7054));
  DFRQX1 \integer_file_reg[9][18] (.C (rc_gclk_199933), .D (n_68), .Q
       (n_7085));
  DFRQX1 \integer_file_reg[9][19] (.C (rc_gclk_199933), .D (n_1598), .Q
       (n_7116));
  DFRQX1 \integer_file_reg[9][1] (.C (rc_gclk_199933), .D (n_24), .Q
       (n_6496));
  DFRQX1 \integer_file_reg[9][20] (.C (rc_gclk_199933), .D (n_1597), .Q
       (n_7147));
  DFRQX1 \integer_file_reg[9][21] (.C (rc_gclk_199933), .D (n_1596), .Q
       (n_7178));
  DFRQX1 \integer_file_reg[9][22] (.C (rc_gclk_199933), .D (n_1595), .Q
       (n_7209));
  DFRQX1 \integer_file_reg[9][23] (.C (rc_gclk_199933), .D (n_1594), .Q
       (n_6279));
  DFRQX1 \integer_file_reg[9][24] (.C (rc_gclk_199933), .D (n_45), .Q
       (n_6310));
  DFRQX1 \integer_file_reg[9][25] (.C (rc_gclk_199933), .D (n_1593), .Q
       (n_6341));
  DFRQX1 \integer_file_reg[9][26] (.C (rc_gclk_199933), .D (n_16), .Q
       (n_6372));
  DFRQX1 \integer_file_reg[9][27] (.C (rc_gclk_199933), .D (n_1592), .Q
       (n_6403));
  DFRQX1 \integer_file_reg[9][28] (.C (rc_gclk_199933), .D (n_1591), .Q
       (n_6434));
  DFRQX1 \integer_file_reg[9][29] (.C (rc_gclk_199933), .D (n_1590), .Q
       (n_6558));
  DFRQX1 \integer_file_reg[9][2] (.C (rc_gclk_199933), .D (n_54), .Q
       (n_6527));
  DFRQX1 \integer_file_reg[9][30] (.C (rc_gclk_199933), .D (n_1589), .Q
       (n_6899));
  DFRQX1 \integer_file_reg[9][31] (.C (rc_gclk_199933), .D (n_1588), .Q
       (n_7240));
  DFRQX1 \integer_file_reg[9][3] (.C (rc_gclk_199933), .D (n_38), .Q
       (n_6589));
  DFRQX1 \integer_file_reg[9][4] (.C (rc_gclk_199933), .D (n_29), .Q
       (n_6620));
  DFRQX1 \integer_file_reg[9][5] (.C (rc_gclk_199933), .D (n_23), .Q
       (n_6651));
  DFRQX1 \integer_file_reg[9][6] (.C (rc_gclk_199933), .D (n_46), .Q
       (n_6682));
  DFRQX1 \integer_file_reg[9][7] (.C (rc_gclk_199933), .D (n_74), .Q
       (n_6713));
  DFRQX1 \integer_file_reg[9][8] (.C (rc_gclk_199933), .D (n_72), .Q
       (n_6744));
  DFRQX1 \integer_file_reg[9][9] (.C (rc_gclk_199933), .D (n_89), .Q
       (n_6775));
  DFRQX1 \prev_instruction_reg[0] (.C (rc_gclk_199999), .D (n_1586), .Q
       (prev_instruction[0]));
  DFRQX1 \prev_instruction_reg[10] (.C (rc_gclk_199999), .D (n_1585),
       .Q (prev_instruction[10]));
  DFRQX1 \prev_instruction_reg[12] (.C (rc_gclk_199999), .D (n_1583),
       .Q (prev_instruction[12]));
  DFRQX1 \prev_instruction_reg[13] (.C (rc_gclk_199999), .D (n_1582),
       .Q (prev_instruction[13]));
  DFRQX1 \prev_instruction_reg[14] (.C (rc_gclk_199999), .D (n_1581),
       .Q (prev_instruction[14]));
  DFRQX1 \prev_instruction_reg[15] (.C (rc_gclk_199999), .D (n_1580),
       .Q (prev_instruction[15]));
  DFRQX1 \prev_instruction_reg[16] (.C (rc_gclk_199999), .D (n_1579),
       .Q (prev_instruction[16]));
  DFRQX1 \prev_instruction_reg[17] (.C (rc_gclk_199999), .D (n_1578),
       .Q (prev_instruction[17]));
  DFRQX1 \prev_instruction_reg[18] (.C (rc_gclk_199999), .D (n_1577),
       .Q (prev_instruction[18]));
  DFRQX1 \prev_instruction_reg[19] (.C (rc_gclk_199999), .D (n_1576),
       .Q (prev_instruction[19]));
  DFRQX1 \prev_instruction_reg[1] (.C (rc_gclk_199999), .D (n_1575), .Q
       (prev_instruction[1]));
  DFRQX1 \prev_instruction_reg[20] (.C (rc_gclk_199999), .D (n_1574),
       .Q (prev_instruction[20]));
  DFRQX1 \prev_instruction_reg[21] (.C (rc_gclk_199999), .D (n_1573),
       .Q (prev_instruction[21]));
  DFRQX1 \prev_instruction_reg[22] (.C (rc_gclk_199999), .D (n_1572),
       .Q (prev_instruction[22]));
  DFRQX1 \prev_instruction_reg[23] (.C (rc_gclk_199999), .D (n_1571),
       .Q (prev_instruction[23]));
  DFRQX1 \prev_instruction_reg[24] (.C (rc_gclk_199999), .D (n_1570),
       .Q (prev_instruction[24]));
  DFRQX1 \prev_instruction_reg[25] (.C (rc_gclk_199999), .D (n_1569),
       .Q (prev_instruction[25]));
  DFRQX1 \prev_instruction_reg[26] (.C (rc_gclk_199999), .D (n_1568),
       .Q (prev_instruction[26]));
  DFRQX1 \prev_instruction_reg[27] (.C (rc_gclk_199999), .D (n_1567),
       .Q (prev_instruction[27]));
  DFRQX1 \prev_instruction_reg[28] (.C (rc_gclk_199999), .D (n_1566),
       .Q (prev_instruction[28]));
  DFRQX1 \prev_instruction_reg[29] (.C (rc_gclk_199999), .D (n_1565),
       .Q (prev_instruction[29]));
  DFRQX1 \prev_instruction_reg[2] (.C (rc_gclk_199999), .D (n_1564), .Q
       (prev_instruction[2]));
  DFRQX1 \prev_instruction_reg[30] (.C (rc_gclk_199999), .D (n_1563),
       .Q (prev_instruction[30]));
  DFRQX1 \prev_instruction_reg[31] (.C (rc_gclk_199999), .D (n_1562),
       .Q (prev_instruction[31]));
  DFRQX1 \prev_instruction_reg[3] (.C (rc_gclk_199999), .D (n_1561), .Q
       (prev_instruction[3]));
  DFRQX1 \prev_instruction_reg[4] (.C (rc_gclk_199999), .D (n_1560), .Q
       (prev_instruction[4]));
  DFRQX1 \prev_instruction_reg[5] (.C (rc_gclk_199999), .D (n_1559), .Q
       (prev_instruction[5]));
  DFRQX1 \prev_instruction_reg[6] (.C (rc_gclk_199999), .D (n_1558), .Q
       (prev_instruction[6]));
  DFRQX1 \prev_instruction_reg[7] (.C (rc_gclk_199999), .D (n_1557), .Q
       (prev_instruction[7]));
  DFRQX1 \prev_instruction_reg[8] (.C (rc_gclk_199999), .D (n_1556), .Q
       (prev_instruction[8]));
  DFRQX1 \prev_instruction_reg[9] (.C (rc_gclk_199999), .D (n_1555), .Q
       (prev_instruction[9]));
  DFRQX1 \program_counter_reg[1] (.C (rc_gclk_199879), .D (n_1475), .Q
       (program_counter[1]));
  NA2I1X1 g92621(.B (n_1454), .AN (n_7304), .Q (n_157));
  NA2I1X1 g92622(.B (n_7275), .AN (n_8078), .Q (n_156));
  NA3I1X1 g92623(.B (n_952), .C (n_953), .AN (n_850), .Q (n_155));
  OR2X1 g92624(.A (n_821), .B (n_820), .Q (n_154));
  NA2I1X2 g92625(.B (n_914), .AN (n_494), .Q (n_153));
  NA2I1X1 g92626(.B (alu_2nd_operand[0]), .AN (n_777), .Q (n_152));
  NA2I1X1 g92627(.B (alu_2nd_operand[3]), .AN (n_408), .Q (n_151));
  NA2I1X1 g92628(.B (alu_2nd_operand[23]), .AN (n_6143), .Q (n_150));
  NA2I1X1 g92629(.B (n_8677), .AN (n_898), .Q (n_149));
  NA2I1X1 g92630(.B (alu_2nd_operand[24]), .AN (n_6145), .Q (n_148));
  AND2X1 g54557(.A (n_8496), .B (n_828), .Q (n_167));
  AND2X1 g54559(.A (n_852), .B (n_8487), .Q (n_160));
  AND2X1 g54561(.A (n_7625), .B (n_181), .Q (n_184));
  AND2X1 g54563(.A (n_7626), .B (n_181), .Q (n_183));
  AND2X1 g54565(.A (n_7630), .B (n_181), .Q (n_182));
  INX1 g54567(.A (n_830), .Q (n_170));
  INX2 g54569(.A (n_361), .Q (n_161));
  OA221X1 g54571(.A (n_631), .B (n_489), .C (n_826), .D (n_687), .E
       (n_488), .Q (n_168));
  INX1 g54577(.A (n_166), .Q (n_162));
  AND2X1 g54579(.A (n_167), .B (n_816), .Q (n_165));
  OA221X1 g54581(.A (n_497), .B (n_166), .C (n_631), .D (n_630), .E
       (n_496), .Q (n_169));
  INX2 g54585(.A (alu_2nd_operand[3]), .Q (n_173));
  OA221X1 g54589(.A (n_686), .B (n_343), .C (n_824), .D (n_733), .E
       (n_342), .Q (n_163));
  OA221X1 g54591(.A (n_794), .B (n_985), .C (n_170), .D (n_589), .E
       (n_588), .Q (n_171));
  AND2X1 g54593(.A (n_8354), .B (n_181), .Q (n_147));
  AND2X1 g54596(.A (n_7395), .B (n_181), .Q (n_146));
  AND2X1 g54597(.A (n_7394), .B (n_181), .Q (n_145));
  AND2X1 g54599(.A (n_7393), .B (n_181), .Q (n_144));
  AND2X1 g54601(.A (n_7392), .B (n_181), .Q (n_143));
  AND2X1 g54602(.A (n_7391), .B (n_181), .Q (n_142));
  AND2X1 g54603(.A (n_8622), .B (n_181), .Q (n_141));
  AND2X1 g54604(.A (n_7389), .B (n_181), .Q (n_140));
  AND2X1 g54606(.A (n_7388), .B (n_181), .Q (n_139));
  AND2X1 g54607(.A (n_7387), .B (n_181), .Q (n_138));
  AND2X1 g54610(.A (n_7386), .B (n_181), .Q (n_137));
  AND2X1 g54612(.A (n_7385), .B (n_181), .Q (n_136));
  AND2X1 g54614(.A (n_7384), .B (n_181), .Q (n_135));
  AND2X1 g54615(.A (n_7383), .B (n_181), .Q (n_134));
  AND2X1 g54617(.A (n_8571), .B (n_181), .Q (n_133));
  AND2X1 g54618(.A (n_7381), .B (n_181), .Q (n_132));
  AND2X1 g54620(.A (n_7380), .B (n_181), .Q (n_131));
  AND2X1 g54623(.A (n_7379), .B (n_181), .Q (n_130));
  AND2X1 g54625(.A (n_7378), .B (n_181), .Q (n_129));
  AND2X1 g54626(.A (n_7377), .B (n_181), .Q (n_128));
  AND2X1 g54627(.A (n_6232), .B (n_181), .Q (n_127));
  AND2X1 g54628(.A (n_6237), .B (n_181), .Q (n_126));
  AND2X1 g54630(.A (n_7398), .B (n_181), .Q (n_125));
  AND2X1 g54631(.A (n_7397), .B (n_181), .Q (n_124));
  AND2X1 g54633(.A (n_7376), .B (n_181), .Q (n_123));
  AND2X1 g54634(.A (n_7635), .B (n_181), .Q (n_122));
  AND2X1 g54635(.A (n_7377), .B (n_181), .Q (n_121));
  AND2X1 g54636(.A (n_7381), .B (n_181), .Q (n_120));
  AND2X1 g54637(.A (n_7383), .B (n_181), .Q (n_119));
  AND2X1 g54638(.A (n_7387), .B (n_181), .Q (n_118));
  AND2X1 g54639(.A (n_7389), .B (n_181), .Q (n_117));
  AND2X1 g54640(.A (n_8622), .B (n_181), .Q (n_116));
  AND2X1 g54641(.A (n_6234), .B (n_181), .Q (n_115));
  NO2X1 g54642(.A (n_1447), .B (n_179), .Q (n_114));
  NO2X1 g54647(.A (n_1165), .B (n_1), .Q (n_113));
  NO2X1 g54661(.A (n_1165), .B (n_179), .Q (n_112));
  NO2X2 g54662(.A (n_1165), .B (n_179), .Q (n_111));
  NO2X1 g54669(.A (n_1165), .B (n_1), .Q (n_110));
  NO2X1 g54670(.A (n_1163), .B (n_1), .Q (n_109));
  NO2X1 g54671(.A (n_1163), .B (n_1), .Q (n_108));
  NO2X1 g54672(.A (n_1163), .B (n_1), .Q (n_107));
  NO2X1 g54673(.A (n_1163), .B (n_1), .Q (n_106));
  NO2X1 g54674(.A (n_1163), .B (n_1), .Q (n_105));
  NO2X2 g54691(.A (n_1162), .B (n_1), .Q (n_104));
  NO2X2 g54701(.A (n_1160), .B (n_1), .Q (n_103));
  NO2X1 g54703(.A (n_1138), .B (n_1), .Q (n_102));
  NO2X1 g54712(.A (n_1137), .B (n_179), .Q (n_101));
  NO2X1 g54724(.A (n_1136), .B (n_179), .Q (n_100));
  NO2X1 g54725(.A (n_1136), .B (n_179), .Q (n_99));
  NO2X1 g54732(.A (n_1160), .B (n_1), .Q (n_98));
  NO2X1 g54736(.A (n_1159), .B (n_180), .Q (n_97));
  NO2X1 g54737(.A (n_1159), .B (n_180), .Q (n_96));
  NO2X1 g54738(.A (n_1159), .B (n_180), .Q (n_95));
  NO2X1 g54739(.A (n_1159), .B (n_180), .Q (n_94));
  NO2X1 g54740(.A (n_1159), .B (n_180), .Q (n_93));
  NO2X1 g54741(.A (n_1159), .B (n_180), .Q (n_92));
  NO2X2 g54744(.A (n_1159), .B (n_180), .Q (n_91));
  NO2X1 g54745(.A (n_1138), .B (n_180), .Q (n_90));
  NO2X2 g54755(.A (n_1136), .B (n_1), .Q (n_89));
  NO2X1 g54756(.A (n_1163), .B (n_1), .Q (n_88));
  NO2X1 g54757(.A (n_1163), .B (n_1), .Q (n_87));
  NO2X1 g54758(.A (n_1163), .B (n_1), .Q (n_86));
  NO2X1 g54759(.A (n_1163), .B (n_1), .Q (n_85));
  NO2X1 g54760(.A (n_1163), .B (n_1), .Q (n_84));
  NO2X1 g54761(.A (n_1163), .B (n_1), .Q (n_83));
  NO2X1 g54779(.A (n_1138), .B (n_1), .Q (n_82));
  NO2X1 g54780(.A (n_1138), .B (n_1), .Q (n_81));
  NO2X1 g54791(.A (n_1137), .B (n_1), .Q (n_80));
  NO2X1 g54798(.A (n_1164), .B (n_1), .Q (n_79));
  NO2X1 g54802(.A (n_1136), .B (n_1), .Q (n_78));
  NO2X1 g54806(.A (n_1164), .B (n_1), .Q (n_77));
  NO2X2 g54814(.A (n_1163), .B (n_179), .Q (n_76));
  NO2X2 g54825(.A (n_1160), .B (n_179), .Q (n_75));
  NO2X1 g54829(.A (n_1138), .B (n_179), .Q (n_74));
  NO2X1 g54833(.A (n_1162), .B (n_1), .Q (n_73));
  NO2X1 g54841(.A (n_1137), .B (n_1), .Q (n_72));
  NO2X1 g54848(.A (n_1162), .B (n_179), .Q (n_71));
  NO2X1 g54862(.A (n_1166), .B (n_1), .Q (n_70));
  NO2X1 g54863(.A (n_1166), .B (n_1), .Q (n_69));
  NO2X1 g54864(.A (n_1158), .B (n_180), .Q (n_68));
  NO2X1 g54865(.A (n_1158), .B (n_180), .Q (n_67));
  NO2X1 g54866(.A (n_1158), .B (n_180), .Q (n_66));
  NO2X1 g54867(.A (n_1158), .B (n_180), .Q (n_65));
  NO2X1 g54868(.A (n_1158), .B (n_180), .Q (n_64));
  NO2X1 g54869(.A (n_1158), .B (n_180), .Q (n_63));
  NO2X1 g54870(.A (n_1158), .B (n_180), .Q (n_62));
  NO2X1 g54871(.A (n_1158), .B (n_180), .Q (n_61));
  NO2X1 g54872(.A (n_1158), .B (n_180), .Q (n_60));
  NO2X1 g54873(.A (n_1158), .B (n_180), .Q (n_59));
  NO2X1 g54874(.A (n_1158), .B (n_180), .Q (n_58));
  NO2X1 g54875(.A (n_1158), .B (n_180), .Q (n_57));
  NO2X1 g54876(.A (n_1158), .B (n_180), .Q (n_56));
  NO2X1 g54878(.A (n_1156), .B (n_180), .Q (n_55));
  NO2X1 g54888(.A (n_1145), .B (n_1), .Q (n_54));
  NO2X1 g54894(.A (n_1142), .B (n_1), .Q (n_53));
  NO2X1 g54895(.A (n_1141), .B (n_179), .Q (n_52));
  NO2X1 g54896(.A (n_1141), .B (n_179), .Q (n_51));
  NO2X1 g54897(.A (n_1141), .B (n_179), .Q (n_50));
  NO2X1 g54898(.A (n_1140), .B (n_1), .Q (n_49));
  NO2X1 g54899(.A (n_1140), .B (n_1), .Q (n_48));
  NO2X1 g54900(.A (n_1140), .B (n_1), .Q (n_47));
  NO2X1 g54911(.A (n_1139), .B (n_1), .Q (n_46));
  NO2X1 g54912(.A (n_1151), .B (n_180), .Q (n_45));
  NO2X1 g54913(.A (n_1151), .B (n_180), .Q (n_44));
  NO2X1 g54914(.A (n_1151), .B (n_180), .Q (n_43));
  NO2X1 g54915(.A (n_1151), .B (n_180), .Q (n_42));
  NO2X1 g54916(.A (n_1151), .B (n_180), .Q (n_41));
  NO2X1 g54917(.A (n_1151), .B (n_180), .Q (n_40));
  NO2X2 g54930(.A (n_1145), .B (n_1), .Q (n_39));
  NO2X2 g54942(.A (n_1142), .B (n_179), .Q (n_38));
  NO2X1 g54950(.A (n_1139), .B (n_179), .Q (n_37));
  NO2X1 g54957(.A (n_1166), .B (n_179), .Q (n_36));
  NO2X1 g54961(.A (n_1141), .B (n_1), .Q (n_35));
  NO2X1 g54962(.A (n_1141), .B (n_1), .Q (n_34));
  NO2X2 g54965(.A (n_1141), .B (n_1), .Q (n_33));
  NO2X1 g54980(.A (n_1140), .B (n_179), .Q (n_32));
  NO2X2 g54981(.A (n_1140), .B (n_179), .Q (n_31));
  NO2X1 g54989(.A (n_1156), .B (n_1), .Q (n_30));
  NO2X1 g55000(.A (n_1141), .B (n_1), .Q (n_29));
  NO2X2 g55001(.A (n_1141), .B (n_1), .Q (n_28));
  NO2X1 g55010(.A (n_1139), .B (n_1), .Q (n_27));
  NO2X1 g55015(.A (n_1156), .B (n_179), .Q (n_26));
  NO2X2 g55025(.A (n_1142), .B (n_1), .Q (n_25));
  NO2X2 g55037(.A (n_1156), .B (n_1), .Q (n_24));
  NO2X1 g55043(.A (n_1140), .B (n_1), .Q (n_23));
  NO2X1 g55047(.A (n_1158), .B (n_179), .Q (n_22));
  NO2X1 g55052(.A (n_1145), .B (n_179), .Q (n_21));
  NO2X1 g55057(.A (n_1166), .B (n_1), .Q (n_20));
  NO2X2 g55067(.A (n_1161), .B (n_1), .Q (n_19));
  NO2X2 g55080(.A (n_1161), .B (n_179), .Q (n_18));
  NO2X1 g55085(.A (n_1161), .B (n_1), .Q (n_17));
  NO2X1 g55086(.A (n_1149), .B (n_180), .Q (n_16));
  NO2X1 g55087(.A (n_1149), .B (n_180), .Q (n_15));
  NO2X1 g55088(.A (n_1149), .B (n_180), .Q (n_14));
  NO2X1 g55089(.A (n_1149), .B (n_180), .Q (n_13));
  NO2X1 g55090(.A (n_1149), .B (n_180), .Q (n_12));
  NO2X1 g55091(.A (n_1149), .B (n_180), .Q (n_11));
  NO2X1 g55092(.A (n_1149), .B (n_180), .Q (n_10));
  NO2X1 g55093(.A (n_1149), .B (n_180), .Q (n_9));
  NO2X1 g55094(.A (n_1149), .B (n_180), .Q (n_8));
  NO2X1 g55095(.A (n_1149), .B (n_180), .Q (n_7));
  NO2X1 g55096(.A (n_1149), .B (n_180), .Q (n_6));
  NO2X1 g55097(.A (n_1149), .B (n_179), .Q (n_5));
  NO2X1 g55098(.A (n_1149), .B (n_179), .Q (n_4));
  NO2X1 g55099(.A (n_1149), .B (n_179), .Q (n_3));
  NO2X1 g55100(.A (n_1149), .B (n_179), .Q (n_2));
  INCX12 g55104(.A (n_181), .Q (n_1));
  INCX12 g55106(.A (n_181), .Q (n_180));
  INX2 g55108(.A (n_164), .Q (n_166));
  EN2X1 add_463_14_g965(.A (add_463_14_n_607), .B (add_463_14_n_817),
       .Q (n_7782));
  EN2X1 add_463_14_g966(.A (add_463_14_n_599), .B (add_463_14_n_845),
       .Q (n_7788));
  EN2X1 add_463_14_g967(.A (add_463_14_n_600), .B (add_463_14_n_847),
       .Q (n_7792));
  EN2X1 add_463_14_g968(.A (add_463_14_n_601), .B (add_463_14_n_880),
       .Q (n_7794));
  EN3X1 add_463_14_g969(.A (add_463_14_n_603), .B (n_6134), .C
       (n_8263), .Q (n_7766));
  EN2X1 add_463_14_g970(.A (add_463_14_n_606), .B (add_463_14_n_855),
       .Q (n_7778));
  EN2X1 add_463_14_g971(.A (add_463_14_n_597), .B (add_463_14_n_866),
       .Q (n_7780));
  EN2X1 add_463_14_g972(.A (add_463_14_n_623), .B (add_463_14_n_814),
       .Q (n_7768));
  EN2X1 add_463_14_g973(.A (add_463_14_n_609), .B (add_463_14_n_811),
       .Q (n_7784));
  EN2X1 add_463_14_g974(.A (add_463_14_n_610), .B (add_463_14_n_843),
       .Q (n_7786));
  EN2X1 add_463_14_g975(.A (add_463_14_n_620), .B (add_463_14_n_826),
       .Q (n_7790));
  EN2X1 add_463_14_g976(.A (add_463_14_n_605), .B (add_463_14_n_810),
       .Q (n_7776));
  EN2X1 add_463_14_g977(.A (add_463_14_n_622), .B (add_463_14_n_823),
       .Q (n_7770));
  EN2X1 add_463_14_g978(.A (add_463_14_n_618), .B (add_463_14_n_813),
       .Q (n_7772));
  EN2X1 add_463_14_g979(.A (add_463_14_n_619), .B (add_463_14_n_804),
       .Q (n_7774));
  MU2IX1 add_463_14_g980(.S (add_463_14_n_864), .IN0
       (add_463_14_n_641), .IN1 (add_463_14_n_640), .Q (n_7796));
  AN21X1 add_463_14_g981(.A (add_463_14_n_640), .B (add_463_14_n_726),
       .C (add_463_14_n_683), .Q (add_463_14_n_597));
  AN21X1 add_463_14_g982(.A (add_463_14_n_640), .B (add_463_14_n_762),
       .C (add_463_14_n_709), .Q (add_463_14_n_599));
  AN21X1 add_463_14_g983(.A (add_463_14_n_640), .B (add_463_14_n_838),
       .C (add_463_14_n_779), .Q (add_463_14_n_600));
  ON21X1 add_463_14_g984(.A (add_463_14_n_641), .B (add_463_14_n_944),
       .C (add_463_14_n_946), .Q (add_463_14_n_601));
  AN31X1 add_463_14_g985(.A (add_463_14_n_722), .B (add_463_14_n_726),
       .C (add_463_14_n_640), .D (add_463_14_n_660), .Q
       (add_463_14_n_603));
  AN31X1 add_463_14_g986(.A (add_463_14_n_802), .B (add_463_14_n_726),
       .C (add_463_14_n_640), .D (add_463_14_n_656), .Q
       (add_463_14_n_605));
  AN31X1 add_463_14_g987(.A (add_463_14_n_972), .B (add_463_14_n_726),
       .C (add_463_14_n_640), .D (add_463_14_n_659), .Q
       (add_463_14_n_606));
  AN31X1 add_463_14_g988(.A (add_463_14_n_756), .B (add_463_14_n_762),
       .C (add_463_14_n_640), .D (add_463_14_n_681), .Q
       (add_463_14_n_607));
  AN31X1 add_463_14_g989(.A (add_463_14_n_799), .B (add_463_14_n_762),
       .C (add_463_14_n_640), .D (add_463_14_n_688), .Q
       (add_463_14_n_609));
  AN31X1 add_463_14_g990(.A (add_463_14_n_968), .B (add_463_14_n_762),
       .C (add_463_14_n_640), .D (add_463_14_n_682), .Q
       (add_463_14_n_610));
  EN2X1 add_463_14_g991(.A (add_463_14_n_639), .B (add_463_14_n_877),
       .Q (n_7810));
  EN2X1 add_463_14_g992(.A (add_463_14_n_628), .B (add_463_14_n_853),
       .Q (n_7802));
  EN2X1 add_463_14_g993(.A (n_8342), .B (add_463_14_n_812), .Q
       (n_7800));
  EN2X1 add_463_14_g994(.A (add_463_14_n_625), .B (add_463_14_n_807),
       .Q (n_7798));
  EN2X1 add_463_14_g995(.A (add_463_14_n_634), .B (add_463_14_n_828),
       .Q (n_7806));
  EN2X1 add_463_14_g996(.A (add_463_14_n_636), .B (add_463_14_n_850),
       .Q (n_7808));
  EN2X1 add_463_14_g997(.A (add_463_14_n_632), .B (add_463_14_n_857),
       .Q (n_7804));
  AN31X1 add_463_14_g998(.A (add_463_14_n_763), .B (add_463_14_n_726),
       .C (add_463_14_n_640), .D (add_463_14_n_664), .Q
       (add_463_14_n_618));
  AN31X1 add_463_14_g999(.A (add_463_14_n_754), .B (add_463_14_n_726),
       .C (add_463_14_n_640), .D (add_463_14_n_666), .Q
       (add_463_14_n_619));
  AN31X1 add_463_14_g1000(.A (add_463_14_n_966), .B (add_463_14_n_838),
       .C (add_463_14_n_640), .D (add_463_14_n_711), .Q
       (add_463_14_n_620));
  AN31X1 add_463_14_g1001(.A (add_463_14_n_721), .B (add_463_14_n_726),
       .C (add_463_14_n_640), .D (add_463_14_n_663), .Q
       (add_463_14_n_622));
  AN31X1 add_463_14_g1002(.A (add_463_14_n_724), .B (add_463_14_n_726),
       .C (add_463_14_n_640), .D (add_463_14_n_662), .Q
       (add_463_14_n_623));
  EN2X1 add_463_14_g1003(.A (add_463_14_n_647), .B (add_463_14_n_868),
       .Q (n_7812));
  ON31X1 add_463_14_g1004(.A (add_463_14_n_757), .B (add_463_14_n_761),
       .C (add_463_14_n_647), .D (add_463_14_n_678), .Q
       (add_463_14_n_625));
  ON21X1 add_463_14_g1007(.A (add_463_14_n_647), .B (add_463_14_n_761),
       .C (n_8594), .Q (add_463_14_n_632));
  AN21X1 add_463_14_g1009(.A (add_463_14_n_646), .B (add_463_14_n_839),
       .C (add_463_14_n_780), .Q (add_463_14_n_636));
  ON21X1 add_463_14_g1010(.A (add_463_14_n_647), .B (add_463_14_n_952),
       .C (add_463_14_n_950), .Q (add_463_14_n_639));
  INX2 add_463_14_g1011(.A (add_463_14_n_640), .Q (add_463_14_n_641));
  NA2X4 add_463_14_g1012(.A (n_8592), .B (add_463_14_n_680), .Q
       (add_463_14_n_640));
  EN2X1 add_463_14_g1014(.A (add_463_14_n_648), .B (add_463_14_n_859),
       .Q (n_7816));
  EN2X1 add_463_14_g1015(.A (add_463_14_n_655), .B (add_463_14_n_872),
       .Q (n_7818));
  EN2X1 add_463_14_g1016(.A (add_463_14_n_653), .B (add_463_14_n_821),
       .Q (n_7814));
  INX1 add_463_14_g1017(.A (add_463_14_n_646), .Q (add_463_14_n_647));
  NA2X4 add_463_14_g1018(.A (add_463_14_n_649), .B (add_463_14_n_717),
       .Q (add_463_14_n_646));
  NO2X1 add_463_14_g1019(.A (add_463_14_n_667), .B (add_463_14_n_781),
       .Q (add_463_14_n_648));
  NA2X2 add_463_14_g1020(.A (add_463_14_n_667), .B (add_463_14_n_797),
       .Q (add_463_14_n_649));
  EN2X0 add_463_14_g1021(.A (add_463_14_n_672), .B (add_463_14_n_862),
       .Q (n_7820));
  EN2X1 add_463_14_g1022(.A (add_463_14_n_673), .B (add_463_14_n_875),
       .Q (n_7822));
  AN31X1 add_463_14_g1023(.A (add_463_14_n_974), .B (add_463_14_n_837),
       .C (add_463_14_n_672), .D (add_463_14_n_714), .Q
       (add_463_14_n_653));
  ON21X1 add_463_14_g1024(.A (n_8593), .B (add_463_14_n_953), .C
       (add_463_14_n_947), .Q (add_463_14_n_655));
  AO21X1 add_463_14_g1025(.A (add_463_14_n_683), .B (add_463_14_n_802),
       .C (add_463_14_n_778), .Q (add_463_14_n_656));
  ON21X1 add_463_14_g1026(.A (add_463_14_n_684), .B (add_463_14_n_971),
       .C (add_463_14_n_906), .Q (add_463_14_n_659));
  ON21X1 add_463_14_g1027(.A (add_463_14_n_684), .B (add_463_14_n_723),
       .C (add_463_14_n_676), .Q (add_463_14_n_660));
  ON21X1 add_463_14_g1028(.A (add_463_14_n_684), .B (add_463_14_n_725),
       .C (add_463_14_n_675), .Q (add_463_14_n_662));
  ON221X1 add_463_14_g1029(.A (add_463_14_n_720), .B
       (add_463_14_n_684), .C (add_463_14_n_917), .D
       (add_463_14_n_697), .E (add_463_14_n_899), .Q
       (add_463_14_n_663));
  ON21X1 add_463_14_g1030(.A (add_463_14_n_684), .B (add_463_14_n_764),
       .C (add_463_14_n_697), .Q (add_463_14_n_664));
  ON211X1 add_463_14_g1031(.A (add_463_14_n_684), .B
       (add_463_14_n_755), .C (add_463_14_n_730), .D
       (add_463_14_n_895), .Q (add_463_14_n_666));
  EN2X1 add_463_14_g1033(.A (add_463_14_n_691), .B (add_463_14_n_870),
       .Q (n_7824));
  INX1 add_463_14_g1034(.A (n_8593), .Q (add_463_14_n_672));
  AN21X1 add_463_14_g1036(.A (add_463_14_n_691), .B (add_463_14_n_951),
       .C (add_463_14_n_949), .Q (add_463_14_n_673));
  AN21X1 add_463_14_g1037(.A (add_463_14_n_698), .B (add_463_14_n_798),
       .C (add_463_14_n_751), .Q (add_463_14_n_675));
  AN21X1 add_463_14_g1038(.A (add_463_14_n_698), .B (add_463_14_n_753),
       .C (add_463_14_n_701), .Q (add_463_14_n_676));
  AN21X1 add_463_14_g1039(.A (add_463_14_n_699), .B (add_463_14_n_758),
       .C (add_463_14_n_702), .Q (add_463_14_n_678));
  AN21X1 add_463_14_g1040(.A (add_463_14_n_699), .B (add_463_14_n_752),
       .C (add_463_14_n_705), .Q (add_463_14_n_680));
  ON211X1 add_463_14_g1041(.A (add_463_14_n_782), .B
       (add_463_14_n_916), .C (add_463_14_n_693), .D
       (add_463_14_n_905), .Q (add_463_14_n_681));
  ON21X1 add_463_14_g1042(.A (add_463_14_n_710), .B (add_463_14_n_967),
       .C (add_463_14_n_896), .Q (add_463_14_n_682));
  INX2 add_463_14_g1043(.A (add_463_14_n_683), .Q (add_463_14_n_684));
  AO21X2 add_463_14_g1044(.A (add_463_14_n_709), .B (add_463_14_n_759),
       .C (add_463_14_n_703), .Q (add_463_14_n_683));
  NA2X1 add_463_14_g1046(.A (add_463_14_n_695), .B (add_463_14_n_782),
       .Q (add_463_14_n_688));
  INX1 add_463_14_g1048(.A (add_463_14_n_708), .Q (add_463_14_n_691));
  NA2X1 add_463_14_g1049(.A (add_463_14_n_709), .B (add_463_14_n_756),
       .Q (add_463_14_n_693));
  NA2X1 add_463_14_g1050(.A (add_463_14_n_709), .B (add_463_14_n_799),
       .Q (add_463_14_n_695));
  INX1 add_463_14_g1051(.A (add_463_14_n_698), .Q (add_463_14_n_697));
  INX1 add_463_14_g1052(.A (n_8594), .Q (add_463_14_n_699));
  ON21X1 add_463_14_g1053(.A (add_463_14_n_750), .B (add_463_14_n_900),
       .C (add_463_14_n_887), .Q (add_463_14_n_701));
  ON21X1 add_463_14_g1054(.A (add_463_14_n_777), .B (add_463_14_n_913),
       .C (add_463_14_n_910), .Q (add_463_14_n_702));
  ON221X1 add_463_14_g1055(.A (add_463_14_n_782), .B
       (add_463_14_n_793), .C (add_463_14_n_905), .D
       (add_463_14_n_909), .E (add_463_14_n_886), .Q
       (add_463_14_n_703));
  ON211X1 add_463_14_g1056(.A (add_463_14_n_898), .B
       (add_463_14_n_910), .C (add_463_14_n_741), .D
       (add_463_14_n_885), .Q (add_463_14_n_705));
  ON211X1 add_463_14_g1057(.A (add_463_14_n_894), .B
       (add_463_14_n_895), .C (add_463_14_n_740), .D
       (add_463_14_n_888), .Q (add_463_14_n_698));
  INX1 add_463_14_g1059(.A (add_463_14_n_709), .Q (add_463_14_n_710));
  AO21X1 add_463_14_g1060(.A (add_463_14_n_779), .B (add_463_14_n_966),
       .C (add_463_14_n_911), .Q (add_463_14_n_711));
  AO21X1 add_463_14_g1061(.A (add_463_14_n_781), .B (add_463_14_n_974),
       .C (add_463_14_n_907), .Q (add_463_14_n_714));
  AN21X1 add_463_14_g1062(.A (add_463_14_n_797), .B (add_463_14_n_781),
       .C (add_463_14_n_785), .Q (add_463_14_n_717));
  NO2X2 add_463_14_g1064(.A (add_463_14_n_746), .B (add_463_14_n_936),
       .Q (add_463_14_n_708));
  AO21X4 add_463_14_g1065(.A (add_463_14_n_796), .B (add_463_14_n_779),
       .C (add_463_14_n_784), .Q (add_463_14_n_709));
  INX1 add_463_14_g1066(.A (add_463_14_n_721), .Q (add_463_14_n_720));
  INX1 add_463_14_g1067(.A (add_463_14_n_723), .Q (add_463_14_n_722));
  INX1 add_463_14_g1068(.A (add_463_14_n_725), .Q (add_463_14_n_724));
  NA2X1 add_463_14_g1069(.A (add_463_14_n_778), .B (add_463_14_n_914),
       .Q (add_463_14_n_730));
  NO2X1 add_463_14_g1071(.A (add_463_14_n_764), .B (add_463_14_n_917),
       .Q (add_463_14_n_721));
  NA2X1 add_463_14_g1072(.A (add_463_14_n_763), .B (add_463_14_n_753),
       .Q (add_463_14_n_723));
  NA2X1 add_463_14_g1073(.A (add_463_14_n_763), .B (add_463_14_n_798),
       .Q (add_463_14_n_725));
  NA2X1 add_463_14_g1075(.A (add_463_14_n_778), .B (add_463_14_n_794),
       .Q (add_463_14_n_740));
  NA2X1 add_463_14_g1076(.A (add_463_14_n_776), .B (add_463_14_n_795),
       .Q (add_463_14_n_741));
  NO2X2 add_463_14_g1080(.A (add_463_14_n_748), .B (add_463_14_n_938),
       .Q (add_463_14_n_746));
  INX1 add_463_14_g1081(.A (add_463_14_n_749), .Q (add_463_14_n_748));
  INX1 add_463_14_g1082(.A (add_463_14_n_751), .Q (add_463_14_n_750));
  INX1 add_463_14_g1083(.A (add_463_14_n_755), .Q (add_463_14_n_754));
  INX1 add_463_14_g1084(.A (add_463_14_n_758), .Q (add_463_14_n_757));
  INX1 add_463_14_g1085(.A (add_463_14_n_760), .Q (add_463_14_n_761));
  INX1 add_463_14_g1086(.A (add_463_14_n_763), .Q (add_463_14_n_764));
  HAX2 add_463_14_g1087(.A (n_6121), .B (n_7692), .S (n_7828), .CO
       (add_463_14_n_749));
  ON21X1 add_463_14_g1088(.A (add_463_14_n_897), .B (add_463_14_n_899),
       .C (add_463_14_n_884), .Q (add_463_14_n_751));
  AND2X1 add_463_14_g1089(.A (add_463_14_n_795), .B (add_463_14_n_800),
       .Q (add_463_14_n_752));
  NO2I1X1 add_463_14_g1090(.B (add_463_14_n_900), .AN
       (add_463_14_n_798), .Q (add_463_14_n_753));
  NA2X1 add_463_14_g1091(.A (add_463_14_n_802), .B (add_463_14_n_914),
       .Q (add_463_14_n_755));
  NO2I1X1 add_463_14_g1092(.B (add_463_14_n_916), .AN
       (add_463_14_n_799), .Q (add_463_14_n_756));
  NO2X1 add_463_14_g1093(.A (add_463_14_n_801), .B (add_463_14_n_913),
       .Q (add_463_14_n_758));
  NO2I1X1 add_463_14_g1094(.B (add_463_14_n_793), .AN
       (add_463_14_n_799), .Q (add_463_14_n_759));
  AND2X2 add_463_14_g1097(.A (add_463_14_n_794), .B (add_463_14_n_802),
       .Q (add_463_14_n_763));
  INX1 add_463_14_g1098(.A (add_463_14_n_776), .Q (add_463_14_n_777));
  ON21X1 add_463_14_g1099(.A (add_463_14_n_955), .B (add_463_14_n_904),
       .C (add_463_14_n_889), .Q (add_463_14_n_783));
  ON21X1 add_463_14_g1100(.A (add_463_14_n_956), .B (add_463_14_n_912),
       .C (add_463_14_n_891), .Q (add_463_14_n_784));
  ON21X1 add_463_14_g1101(.A (add_463_14_n_954), .B (add_463_14_n_908),
       .C (add_463_14_n_893), .Q (add_463_14_n_785));
  ON21X1 add_463_14_g1103(.A (add_463_14_n_962), .B (add_463_14_n_901),
       .C (add_463_14_n_883), .Q (add_463_14_n_776));
  ON21X1 add_463_14_g1104(.A (add_463_14_n_945), .B (add_463_14_n_906),
       .C (add_463_14_n_890), .Q (add_463_14_n_778));
  ON21X1 add_463_14_g1105(.A (add_463_14_n_946), .B (add_463_14_n_961),
       .C (add_463_14_n_940), .Q (add_463_14_n_779));
  ON21X1 add_463_14_g1106(.A (add_463_14_n_950), .B (add_463_14_n_959),
       .C (add_463_14_n_942), .Q (add_463_14_n_780));
  ON21X1 add_463_14_g1107(.A (add_463_14_n_947), .B (add_463_14_n_960),
       .C (add_463_14_n_941), .Q (add_463_14_n_781));
  OA21X2 add_463_14_g1108(.A (add_463_14_n_957), .B (add_463_14_n_896),
       .C (add_463_14_n_892), .Q (add_463_14_n_782));
  INX1 add_463_14_g1109(.A (add_463_14_n_800), .Q (add_463_14_n_801));
  NO2X1 add_463_14_g1110(.A (add_463_14_n_955), .B (add_463_14_n_969),
       .Q (add_463_14_n_792));
  NO2I1X1 add_463_14_g1111(.B (add_463_14_n_894), .AN
       (add_463_14_n_888), .Q (add_463_14_n_804));
  NA2I1X1 add_463_14_g1112(.B (add_463_14_n_885), .AN
       (add_463_14_n_898), .Q (add_463_14_n_807));
  AND2X1 add_463_14_g1113(.A (add_463_14_n_914), .B (add_463_14_n_895),
       .Q (add_463_14_n_810));
  NO2I1X1 add_463_14_g1114(.B (add_463_14_n_916), .AN
       (add_463_14_n_905), .Q (add_463_14_n_811));
  NO2I1X1 add_463_14_g1115(.B (add_463_14_n_913), .AN
       (add_463_14_n_910), .Q (add_463_14_n_812));
  NO2I1X1 add_463_14_g1116(.B (add_463_14_n_917), .AN
       (add_463_14_n_899), .Q (add_463_14_n_813));
  NO2I1X1 add_463_14_g1117(.B (add_463_14_n_900), .AN
       (add_463_14_n_887), .Q (add_463_14_n_814));
  OR2X1 add_463_14_g1118(.A (add_463_14_n_909), .B (add_463_14_n_916),
       .Q (add_463_14_n_793));
  NO2X1 add_463_14_g1119(.A (add_463_14_n_894), .B (add_463_14_n_915),
       .Q (add_463_14_n_794));
  NO2X1 add_463_14_g1120(.A (add_463_14_n_898), .B (add_463_14_n_913),
       .Q (add_463_14_n_795));
  NO2I1X1 add_463_14_g1121(.B (add_463_14_n_909), .AN
       (add_463_14_n_886), .Q (add_463_14_n_817));
  NO2X1 add_463_14_g1122(.A (add_463_14_n_956), .B (add_463_14_n_965),
       .Q (add_463_14_n_796));
  NO2X1 add_463_14_g1123(.A (add_463_14_n_954), .B (add_463_14_n_973),
       .Q (add_463_14_n_797));
  NO2I1X1 add_463_14_g1124(.B (add_463_14_n_954), .AN
       (add_463_14_n_893), .Q (add_463_14_n_821));
  NO2I1X1 add_463_14_g1125(.B (add_463_14_n_897), .AN
       (add_463_14_n_884), .Q (add_463_14_n_823));
  NO2I1X1 add_463_14_g1126(.B (add_463_14_n_956), .AN
       (add_463_14_n_891), .Q (add_463_14_n_826));
  NA2I1X1 add_463_14_g1127(.B (add_463_14_n_889), .AN
       (add_463_14_n_955), .Q (add_463_14_n_828));
  NO2X1 add_463_14_g1128(.A (add_463_14_n_917), .B (add_463_14_n_897),
       .Q (add_463_14_n_798));
  NO2X1 add_463_14_g1129(.A (add_463_14_n_967), .B (add_463_14_n_957),
       .Q (add_463_14_n_799));
  NO2X1 add_463_14_g1130(.A (add_463_14_n_964), .B (add_463_14_n_962),
       .Q (add_463_14_n_800));
  NO2X1 add_463_14_g1131(.A (add_463_14_n_971), .B (add_463_14_n_945),
       .Q (add_463_14_n_802));
  NA2I1X1 add_463_14_g1133(.B (add_463_14_n_951), .AN
       (add_463_14_n_958), .Q (add_463_14_n_840));
  NO2I1X1 add_463_14_g1134(.B (add_463_14_n_957), .AN
       (add_463_14_n_892), .Q (add_463_14_n_843));
  AND2X1 add_463_14_g1135(.A (add_463_14_n_968), .B (add_463_14_n_896),
       .Q (add_463_14_n_845));
  NO2X1 add_463_14_g1136(.A (add_463_14_n_911), .B (add_463_14_n_965),
       .Q (add_463_14_n_847));
  NO2X1 add_463_14_g1137(.A (add_463_14_n_903), .B (add_463_14_n_969),
       .Q (add_463_14_n_850));
  NA2I1X1 add_463_14_g1138(.B (add_463_14_n_883), .AN
       (add_463_14_n_962), .Q (add_463_14_n_853));
  NO2I1X1 add_463_14_g1139(.B (add_463_14_n_945), .AN
       (add_463_14_n_890), .Q (add_463_14_n_855));
  NA2X1 add_463_14_g1140(.A (add_463_14_n_963), .B (add_463_14_n_901),
       .Q (add_463_14_n_857));
  NO2X1 add_463_14_g1141(.A (add_463_14_n_907), .B (add_463_14_n_973),
       .Q (add_463_14_n_859));
  NA2I1X1 add_463_14_g1142(.B (add_463_14_n_947), .AN
       (add_463_14_n_953), .Q (add_463_14_n_862));
  NO2I1X1 add_463_14_g1143(.B (add_463_14_n_944), .AN
       (add_463_14_n_946), .Q (add_463_14_n_864));
  AND2X1 add_463_14_g1144(.A (add_463_14_n_972), .B (add_463_14_n_906),
       .Q (add_463_14_n_866));
  NO2I1X1 add_463_14_g1145(.B (add_463_14_n_952), .AN
       (add_463_14_n_950), .Q (add_463_14_n_868));
  NA2X1 add_463_14_g1146(.A (add_463_14_n_951), .B (add_463_14_n_948),
       .Q (add_463_14_n_870));
  NA2X1 add_463_14_g1147(.A (add_463_14_n_1078), .B (add_463_14_n_937),
       .Q (add_463_14_n_836));
  NA2I1X1 add_463_14_g1148(.B (add_463_14_n_941), .AN
       (add_463_14_n_960), .Q (add_463_14_n_872));
  NO2X1 add_463_14_g1149(.A (add_463_14_n_953), .B (add_463_14_n_960),
       .Q (add_463_14_n_837));
  NO2I1X1 add_463_14_g1150(.B (add_463_14_n_958), .AN
       (add_463_14_n_943), .Q (add_463_14_n_875));
  NA2I1X1 add_463_14_g1151(.B (add_463_14_n_942), .AN
       (add_463_14_n_959), .Q (add_463_14_n_877));
  NA2I1X1 add_463_14_g1152(.B (add_463_14_n_940), .AN
       (add_463_14_n_961), .Q (add_463_14_n_880));
  NO2X1 add_463_14_g1153(.A (add_463_14_n_944), .B (add_463_14_n_961),
       .Q (add_463_14_n_838));
  NO2X1 add_463_14_g1154(.A (add_463_14_n_952), .B (add_463_14_n_959),
       .Q (add_463_14_n_839));
  INX1 add_463_14_g1155(.A (add_463_14_n_901), .Q (add_463_14_n_902));
  INX1 add_463_14_g1156(.A (add_463_14_n_904), .Q (add_463_14_n_903));
  INX1 add_463_14_g1157(.A (add_463_14_n_908), .Q (add_463_14_n_907));
  INX1 add_463_14_g1158(.A (add_463_14_n_912), .Q (add_463_14_n_911));
  INX1 add_463_14_g1159(.A (add_463_14_n_915), .Q (add_463_14_n_914));
  NA2X1 add_463_14_g1160(.A (\rs1_data[13]_39536 ), .B (n_7689), .Q
       (add_463_14_n_883));
  NA2X1 add_463_14_g1161(.A (\rs1_data[29]_39416 ), .B (n_7672), .Q
       (add_463_14_n_884));
  NA2X1 add_463_14_g1162(.A (\rs1_data[15]_39556 ), .B (n_7687), .Q
       (add_463_14_n_885));
  NA2X1 add_463_14_g1163(.A (\rs1_data[23]_39326 ), .B (n_7678), .Q
       (add_463_14_n_886));
  NA2X1 add_463_14_g1164(.A (\rs1_data[30]_39526 ), .B (n_7671), .Q
       (add_463_14_n_887));
  NA2X1 add_463_14_g1165(.A (n_6135), .B (n_7674), .Q
       (add_463_14_n_888));
  NA2X1 add_463_14_g1166(.A (\rs1_data[11]_39506 ), .B (n_7691), .Q
       (add_463_14_n_889));
  NA2X1 add_463_14_g1167(.A (\rs1_data[25]_39346 ), .B (n_7676), .Q
       (add_463_14_n_890));
  NA2X1 add_463_14_g1168(.A (\rs1_data[19]_39596 ), .B (n_7683), .Q
       (add_463_14_n_891));
  NA2X1 add_463_14_g1169(.A (\rs1_data[21]_39616 ), .B (n_7693), .Q
       (add_463_14_n_892));
  NA2X1 add_463_14_g1170(.A (\rs1_data[7]_39466 ), .B (n_8259), .Q
       (add_463_14_n_893));
  NO2X1 add_463_14_g1171(.A (n_6135), .B (n_7674), .Q
       (add_463_14_n_894));
  NA2X1 add_463_14_g1172(.A (\rs1_data[26]_39356 ), .B (n_7675), .Q
       (add_463_14_n_895));
  NA2X1 add_463_14_g1173(.A (n_6149), .B (n_7670), .Q
       (add_463_14_n_896));
  NO2X1 add_463_14_g1174(.A (\rs1_data[29]_39416 ), .B (n_7672), .Q
       (add_463_14_n_897));
  NO2X1 add_463_14_g1175(.A (\rs1_data[15]_39556 ), .B (n_7687), .Q
       (add_463_14_n_898));
  NA2X1 add_463_14_g1176(.A (n_6136), .B (n_7673), .Q
       (add_463_14_n_899));
  NO2X1 add_463_14_g1177(.A (\rs1_data[30]_39526 ), .B (n_7671), .Q
       (add_463_14_n_900));
  NA2X1 add_463_14_g1178(.A (\rs1_data[12]_39516 ), .B (n_7690), .Q
       (add_463_14_n_901));
  NA2X1 add_463_14_g1179(.A (\rs1_data[10]_39496 ), .B (n_8262), .Q
       (add_463_14_n_904));
  NA2X1 add_463_14_g1180(.A (\rs1_data[22]_39626 ), .B (n_7669), .Q
       (add_463_14_n_905));
  NA2X1 add_463_14_g1181(.A (\rs1_data[24]_39336 ), .B (n_7677), .Q
       (add_463_14_n_906));
  NA2X1 add_463_14_g1182(.A (n_6126), .B (n_8258), .Q
       (add_463_14_n_908));
  NO2X1 add_463_14_g1183(.A (\rs1_data[23]_39326 ), .B (n_7678), .Q
       (add_463_14_n_909));
  NA2X1 add_463_14_g1184(.A (\rs1_data[14]_39546 ), .B (n_7688), .Q
       (add_463_14_n_910));
  NA2X1 add_463_14_g1185(.A (n_6141), .B (n_7684), .Q
       (add_463_14_n_912));
  NO2X1 add_463_14_g1186(.A (\rs1_data[14]_39546 ), .B (n_7688), .Q
       (add_463_14_n_913));
  NO2X1 add_463_14_g1187(.A (\rs1_data[26]_39356 ), .B (n_7675), .Q
       (add_463_14_n_915));
  NO2X1 add_463_14_g1188(.A (\rs1_data[22]_39626 ), .B (n_7669), .Q
       (add_463_14_n_916));
  NO2X1 add_463_14_g1189(.A (n_6136), .B (n_7673), .Q
       (add_463_14_n_917));
  INX1 add_463_14_g1190(.A (add_463_14_n_937), .Q (add_463_14_n_936));
  INX1 add_463_14_g1191(.A (add_463_14_n_1078), .Q (add_463_14_n_938));
  INX1 add_463_14_g1192(.A (add_463_14_n_948), .Q (add_463_14_n_949));
  INX1 add_463_14_g1193(.A (add_463_14_n_964), .Q (add_463_14_n_963));
  INX1 add_463_14_g1194(.A (add_463_14_n_965), .Q (add_463_14_n_966));
  INX1 add_463_14_g1195(.A (add_463_14_n_967), .Q (add_463_14_n_968));
  INX1 add_463_14_g1196(.A (add_463_14_n_969), .Q (add_463_14_n_970));
  INX1 add_463_14_g1197(.A (add_463_14_n_971), .Q (add_463_14_n_972));
  INX1 add_463_14_g1198(.A (add_463_14_n_973), .Q (add_463_14_n_974));
  NA2X1 add_463_14_g1199(.A (\rs1_data[1]_39396 ), .B (n_7682), .Q
       (add_463_14_n_937));
  NA2X1 add_463_14_g1201(.A (n_8366), .B (n_7685), .Q
       (add_463_14_n_940));
  NA2X1 add_463_14_g1202(.A (n_2306), .B (n_8257), .Q
       (add_463_14_n_941));
  NA2X1 add_463_14_g1203(.A (\rs1_data[9]_39486 ), .B (n_8261), .Q
       (add_463_14_n_942));
  NA2X1 add_463_14_g1204(.A (\rs1_data[3]_39426 ), .B (n_7680), .Q
       (add_463_14_n_943));
  NO2X1 add_463_14_g1205(.A (n_6132), .B (n_7686), .Q
       (add_463_14_n_944));
  NO2X1 add_463_14_g1206(.A (\rs1_data[25]_39346 ), .B (n_7676), .Q
       (add_463_14_n_945));
  NA2X1 add_463_14_g1207(.A (n_6132), .B (n_7686), .Q
       (add_463_14_n_946));
  NA2X1 add_463_14_g1208(.A (\rs1_data[4]_39436 ), .B (n_2437), .Q
       (add_463_14_n_947));
  NA2X1 add_463_14_g1209(.A (n_6123), .B (n_7681), .Q
       (add_463_14_n_948));
  NA2X1 add_463_14_g1210(.A (n_6127), .B (n_8260), .Q
       (add_463_14_n_950));
  OR2X1 add_463_14_g1211(.A (n_6123), .B (n_7681), .Q
       (add_463_14_n_951));
  NO2X1 add_463_14_g1212(.A (n_6127), .B (n_8260), .Q
       (add_463_14_n_952));
  NO2X1 add_463_14_g1213(.A (\rs1_data[4]_39436 ), .B (n_2437), .Q
       (add_463_14_n_953));
  NO2X1 add_463_14_g1214(.A (\rs1_data[7]_39466 ), .B (n_8259), .Q
       (add_463_14_n_954));
  NO2X1 add_463_14_g1215(.A (\rs1_data[11]_39506 ), .B (n_7691), .Q
       (add_463_14_n_955));
  NO2X1 add_463_14_g1216(.A (\rs1_data[19]_39596 ), .B (n_7683), .Q
       (add_463_14_n_956));
  NO2X1 add_463_14_g1217(.A (\rs1_data[21]_39616 ), .B (n_7693), .Q
       (add_463_14_n_957));
  NO2X1 add_463_14_g1218(.A (\rs1_data[3]_39426 ), .B (n_7680), .Q
       (add_463_14_n_958));
  NO2X1 add_463_14_g1219(.A (\rs1_data[9]_39486 ), .B (n_8261), .Q
       (add_463_14_n_959));
  NO2X1 add_463_14_g1220(.A (n_2306), .B (n_8257), .Q
       (add_463_14_n_960));
  NO2X1 add_463_14_g1221(.A (n_8366), .B (n_7685), .Q
       (add_463_14_n_961));
  NO2X1 add_463_14_g1222(.A (\rs1_data[13]_39536 ), .B (n_7689), .Q
       (add_463_14_n_962));
  NO2X1 add_463_14_g1223(.A (\rs1_data[12]_39516 ), .B (n_7690), .Q
       (add_463_14_n_964));
  NO2X1 add_463_14_g1224(.A (n_6141), .B (n_7684), .Q
       (add_463_14_n_965));
  NO2X1 add_463_14_g1225(.A (n_6149), .B (n_7670), .Q
       (add_463_14_n_967));
  NO2X1 add_463_14_g1226(.A (\rs1_data[10]_39496 ), .B (n_8262), .Q
       (add_463_14_n_969));
  NO2X1 add_463_14_g1227(.A (\rs1_data[24]_39336 ), .B (n_7677), .Q
       (add_463_14_n_971));
  NO2X1 add_463_14_g1228(.A (n_6126), .B (n_8258), .Q
       (add_463_14_n_973));
  OR2X2 add_463_14_g1231(.A (\rs1_data[1]_39396 ), .B (n_7682), .Q
       (add_463_14_n_1078));
  AND2X1 add_463_14_g1233(.A (add_463_14_n_796), .B (add_463_14_n_838),
       .Q (add_463_14_n_762));
  AO321X1 add_463_14_g1235(.A (add_463_14_n_963), .B
       (add_463_14_n_760), .C (add_463_14_n_646), .D
       (add_463_14_n_963), .E (add_463_14_n_699), .F
       (add_463_14_n_902), .Q (add_463_14_n_628));
  AO321X1 add_463_14_g1237(.A (add_463_14_n_970), .B
       (add_463_14_n_839), .C (add_463_14_n_646), .D
       (add_463_14_n_970), .E (add_463_14_n_780), .F
       (add_463_14_n_903), .Q (add_463_14_n_634));
  NO2I1X2 add_463_14_g1239(.B (n_8593), .AN (add_463_14_n_837), .Q
       (add_463_14_n_667));
  AND2X1 add_463_14_g1241(.A (add_463_14_n_792), .B (add_463_14_n_839),
       .Q (add_463_14_n_760));
  EN2X1 add_464_21_g962(.A (add_464_21_n_596), .B (add_464_21_n_827),
       .Q (n_7779));
  EN2X1 add_464_21_g963(.A (add_464_21_n_626), .B (add_464_21_n_798),
       .Q (n_7767));
  EN2X1 add_464_21_g964(.A (add_464_21_n_625), .B (add_464_21_n_772),
       .Q (n_7769));
  EN2X1 add_464_21_g965(.A (add_464_21_n_622), .B (add_464_21_n_815),
       .Q (n_7773));
  EN2X1 add_464_21_g966(.A (n_8344), .B (add_464_21_n_821), .Q
       (n_7775));
  EN2X1 add_464_21_g967(.A (add_464_21_n_605), .B (add_464_21_n_835),
       .Q (n_7777));
  EN2X1 add_464_21_g969(.A (n_8348), .B (add_464_21_n_779), .Q
       (n_7789));
  EN2X1 add_464_21_g970(.A (n_8346), .B (add_464_21_n_823), .Q
       (n_7783));
  EN2X1 add_464_21_g971(.A (add_464_21_n_611), .B (add_464_21_n_832),
       .Q (n_7785));
  EN2X1 add_464_21_g972(.A (add_464_21_n_597), .B (add_464_21_n_825),
       .Q (n_7787));
  EN2X1 add_464_21_g973(.A (add_464_21_n_608), .B (add_464_21_n_818),
       .Q (n_7781));
  EN2X1 add_464_21_g974(.A (add_464_21_n_599), .B (add_464_21_n_790),
       .Q (n_7791));
  EN2X1 add_464_21_g975(.A (add_464_21_n_600), .B (add_464_21_n_795),
       .Q (n_7793));
  EN2X1 add_464_21_g976(.A (add_464_21_n_621), .B (add_464_21_n_829),
       .Q (n_7771));
  EN2X0 add_464_21_g977(.A (add_464_21_n_638), .B (add_464_21_n_791),
       .Q (n_7795));
  AN21X1 add_464_21_g978(.A (add_464_21_n_637), .B (add_464_21_n_708),
       .C (add_464_21_n_686), .Q (add_464_21_n_596));
  AN21X1 add_464_21_g979(.A (add_464_21_n_637), .B (add_464_21_n_730),
       .C (add_464_21_n_701), .Q (add_464_21_n_597));
  AN21X1 add_464_21_g980(.A (add_464_21_n_637), .B (add_464_21_n_768),
       .C (add_464_21_n_729), .Q (add_464_21_n_599));
  ON21X1 add_464_21_g981(.A (add_464_21_n_638), .B (add_464_21_n_870),
       .C (add_464_21_n_860), .Q (add_464_21_n_600));
  AN31X1 add_464_21_g982(.A (add_464_21_n_714), .B (add_464_21_n_708),
       .C (add_464_21_n_637), .D (add_464_21_n_665), .Q
       (add_464_21_n_602));
  AN31X1 add_464_21_g985(.A (add_464_21_n_745), .B (add_464_21_n_730),
       .C (add_464_21_n_637), .D (add_464_21_n_680), .Q
       (add_464_21_n_608));
  EN2X1 add_464_21_g988(.A (add_464_21_n_632), .B (add_464_21_n_793),
       .Q (n_7799));
  EN2X0 add_464_21_g989(.A (add_464_21_n_648), .B (add_464_21_n_841),
       .Q (n_7809));
  EN2X1 add_464_21_g990(.A (add_464_21_n_645), .B (add_464_21_n_830),
       .Q (n_7807));
  EN2X1 add_464_21_g991(.A (add_464_21_n_643), .B (add_464_21_n_804),
       .Q (n_7805));
  EN2X1 add_464_21_g992(.A (add_464_21_n_642), .B (add_464_21_n_788),
       .Q (n_7803));
  EN2X1 add_464_21_g993(.A (add_464_21_n_634), .B (add_464_21_n_785),
       .Q (n_7797));
  EN2X1 add_464_21_g994(.A (add_464_21_n_639), .B (add_464_21_n_801),
       .Q (n_7801));
  AN31X1 add_464_21_g995(.A (add_464_21_n_754), .B (add_464_21_n_708),
       .C (add_464_21_n_637), .D (add_464_21_n_664), .Q
       (add_464_21_n_621));
  AN31X1 add_464_21_g996(.A (add_464_21_n_749), .B (add_464_21_n_708),
       .C (add_464_21_n_637), .D (n_8595), .Q (add_464_21_n_622));
  AN31X1 add_464_21_g998(.A (add_464_21_n_721), .B (add_464_21_n_708),
       .C (add_464_21_n_637), .D (add_464_21_n_669), .Q
       (add_464_21_n_625));
  NA2X1 add_464_21_g999(.A (add_464_21_n_627), .B (add_464_21_n_667),
       .Q (add_464_21_n_626));
  NA3X1 add_464_21_g1000(.A (add_464_21_n_637), .B (add_464_21_n_708),
       .C (add_464_21_n_717), .Q (add_464_21_n_627));
  EN2X1 add_464_21_g1001(.A (add_464_21_n_654), .B (add_464_21_n_846),
       .Q (n_7811));
  EN2X0 add_464_21_g1002(.A (add_464_21_n_657), .B (add_464_21_n_838),
       .Q (n_7813));
  EN2X0 add_464_21_g1003(.A (add_464_21_n_655), .B (add_464_21_n_813),
       .Q (n_7815));
  EN2X1 add_464_21_g1004(.A (add_464_21_n_661), .B (add_464_21_n_844),
       .Q (n_7817));
  AN321X1 add_464_21_g1005(.A (add_464_21_n_771), .B
       (add_464_21_n_731), .C (add_464_21_n_653), .D
       (add_464_21_n_771), .E (add_464_21_n_702), .F
       (add_464_21_n_727), .Q (add_464_21_n_632));
  AN31X1 add_464_21_g1006(.A (add_464_21_n_731), .B (add_464_21_n_726),
       .C (add_464_21_n_653), .D (add_464_21_n_687), .Q
       (add_464_21_n_634));
  INX1 add_464_21_g1007(.A (add_464_21_n_637), .Q (add_464_21_n_638));
  AO21X1 add_464_21_g1009(.A (add_464_21_n_653), .B (add_464_21_n_731),
       .C (add_464_21_n_702), .Q (add_464_21_n_642));
  AN21X1 add_464_21_g1011(.A (add_464_21_n_653), .B (add_464_21_n_810),
       .C (add_464_21_n_751), .Q (add_464_21_n_645));
  ON21X1 add_464_21_g1012(.A (add_464_21_n_654), .B (add_464_21_n_937),
       .C (add_464_21_n_928), .Q (add_464_21_n_648));
  AO321X4 add_464_21_g1013(.A (add_464_21_n_731), .B
       (add_464_21_n_725), .C (add_464_21_n_653), .D
       (add_464_21_n_725), .E (add_464_21_n_702), .F
       (add_464_21_n_697), .Q (add_464_21_n_637));
  EN2X0 add_464_21_g1014(.A (add_464_21_n_678), .B (add_464_21_n_777),
       .Q (n_7819));
  EN2X0 add_464_21_g1015(.A (add_464_21_n_676), .B (add_464_21_n_782),
       .Q (n_7821));
  INX1 add_464_21_g1016(.A (add_464_21_n_653), .Q (add_464_21_n_654));
  NA2X4 add_464_21_g1017(.A (add_464_21_n_674), .B (add_464_21_n_695),
       .Q (add_464_21_n_653));
  AN21X1 add_464_21_g1018(.A (add_464_21_n_678), .B (add_464_21_n_770),
       .C (add_464_21_n_728), .Q (add_464_21_n_655));
  AN321X1 add_464_21_g1019(.A (add_464_21_n_948), .B
       (add_464_21_n_770), .C (add_464_21_n_678), .D
       (add_464_21_n_948), .E (add_464_21_n_728), .F
       (add_464_21_n_934), .Q (add_464_21_n_657));
  ON21X1 add_464_21_g1020(.A (add_464_21_n_679), .B (add_464_21_n_864),
       .C (add_464_21_n_876), .Q (add_464_21_n_661));
  ON21X1 add_464_21_g1022(.A (add_464_21_n_685), .B (add_464_21_n_753),
       .C (add_464_21_n_703), .Q (add_464_21_n_664));
  AO21X1 add_464_21_g1023(.A (add_464_21_n_686), .B (add_464_21_n_714),
       .C (add_464_21_n_690), .Q (add_464_21_n_665));
  AN221X1 add_464_21_g1024(.A (add_464_21_n_769), .B
       (add_464_21_n_704), .C (add_464_21_n_717), .D
       (add_464_21_n_686), .E (add_464_21_n_746), .Q
       (add_464_21_n_667));
  ON221X1 add_464_21_g1025(.A (add_464_21_n_720), .B
       (add_464_21_n_685), .C (add_464_21_n_943), .D
       (add_464_21_n_703), .E (add_464_21_n_872), .Q
       (add_464_21_n_669));
  NA3X2 add_464_21_g1027(.A (add_464_21_n_678), .B (add_464_21_n_770),
       .C (add_464_21_n_809), .Q (add_464_21_n_674));
  EN2X0 add_464_21_g1028(.A (add_464_21_n_693), .B (add_464_21_n_775),
       .Q (n_7823));
  AN21X1 add_464_21_g1029(.A (add_464_21_n_693), .B (add_464_21_n_865),
       .C (add_464_21_n_862), .Q (add_464_21_n_676));
  INX1 add_464_21_g1030(.A (add_464_21_n_678), .Q (add_464_21_n_679));
  NA2I1X4 add_464_21_g1031(.B (add_464_21_n_691), .AN
       (add_464_21_n_738), .Q (add_464_21_n_678));
  AO221X1 add_464_21_g1032(.A (add_464_21_n_745), .B
       (add_464_21_n_701), .C (add_464_21_n_750), .D
       (add_464_21_n_939), .E (add_464_21_n_932), .Q
       (add_464_21_n_680));
  INX1 add_464_21_g1034(.A (add_464_21_n_685), .Q (add_464_21_n_686));
  AN21X1 add_464_21_g1035(.A (add_464_21_n_701), .B (add_464_21_n_748),
       .C (add_464_21_n_706), .Q (add_464_21_n_685));
  AO221X1 add_464_21_g1036(.A (add_464_21_n_726), .B
       (add_464_21_n_702), .C (add_464_21_n_727), .D
       (add_464_21_n_879), .E (add_464_21_n_859), .Q
       (add_464_21_n_687));
  ON211X1 add_464_21_g1037(.A (add_464_21_n_703), .B
       (add_464_21_n_747), .C (add_464_21_n_723), .D
       (add_464_21_n_855), .Q (add_464_21_n_690));
  NA3X2 add_464_21_g1038(.A (add_464_21_n_693), .B (add_464_21_n_868),
       .C (add_464_21_n_865), .Q (add_464_21_n_691));
  FAX1 add_464_21_g1039(.A (program_counter[1]), .B (n_7682), .CI
       (add_464_21_n_733), .S (n_7825), .CO (add_464_21_n_693));
  AN21X1 add_464_21_g1040(.A (add_464_21_n_728), .B (add_464_21_n_809),
       .C (add_464_21_n_756), .Q (add_464_21_n_695));
  AO21X1 add_464_21_g1041(.A (add_464_21_n_727), .B (add_464_21_n_766),
       .C (add_464_21_n_737), .Q (add_464_21_n_697));
  NA2X2 add_464_21_g1043(.A (add_464_21_n_713), .B (add_464_21_n_734),
       .Q (add_464_21_n_701));
  AO21X1 add_464_21_g1044(.A (add_464_21_n_767), .B (add_464_21_n_751),
       .C (add_464_21_n_736), .Q (add_464_21_n_702));
  INX1 add_464_21_g1045(.A (add_464_21_n_703), .Q (add_464_21_n_704));
  AN21X1 add_464_21_g1046(.A (add_464_21_n_752), .B (add_464_21_n_808),
       .C (add_464_21_n_757), .Q (add_464_21_n_703));
  AO21X1 add_464_21_g1047(.A (add_464_21_n_750), .B (add_464_21_n_807),
       .C (add_464_21_n_755), .Q (add_464_21_n_706));
  NA2X1 add_464_21_g1050(.A (add_464_21_n_729), .B (add_464_21_n_765),
       .Q (add_464_21_n_713));
  NO2X1 add_464_21_g1051(.A (add_464_21_n_753), .B (add_464_21_n_747),
       .Q (add_464_21_n_714));
  AND2X1 add_464_21_g1052(.A (add_464_21_n_754), .B (add_464_21_n_769),
       .Q (add_464_21_n_717));
  INX1 add_464_21_g1053(.A (add_464_21_n_721), .Q (add_464_21_n_720));
  NO2X1 add_464_21_g1054(.A (add_464_21_n_753), .B (add_464_21_n_943),
       .Q (add_464_21_n_721));
  NA2X1 add_464_21_g1055(.A (add_464_21_n_746), .B (add_464_21_n_877),
       .Q (add_464_21_n_723));
  HAX2 add_464_21_g1056(.A (n_7692), .B (program_counter[0]), .S
       (n_7827), .CO (add_464_21_n_733));
  AN21X1 add_464_21_g1057(.A (add_464_21_n_871), .B (add_464_21_n_863),
       .C (add_464_21_n_850), .Q (add_464_21_n_734));
  ON21X1 add_464_21_g1058(.A (add_464_21_n_875), .B (add_464_21_n_925),
       .C (add_464_21_n_854), .Q (add_464_21_n_736));
  ON21X1 add_464_21_g1059(.A (add_464_21_n_873), .B (add_464_21_n_858),
       .C (add_464_21_n_851), .Q (add_464_21_n_737));
  ON21X1 add_464_21_g1060(.A (add_464_21_n_869), .B (add_464_21_n_861),
       .C (add_464_21_n_848), .Q (add_464_21_n_738));
  AND2X1 add_464_21_g1061(.A (add_464_21_n_766), .B (add_464_21_n_771),
       .Q (add_464_21_n_725));
  AND2X1 add_464_21_g1062(.A (add_464_21_n_771), .B (add_464_21_n_879),
       .Q (add_464_21_n_726));
  ON21X1 add_464_21_g1063(.A (add_464_21_n_866), .B (add_464_21_n_856),
       .C (add_464_21_n_849), .Q (add_464_21_n_727));
  ON21X1 add_464_21_g1064(.A (add_464_21_n_876), .B (add_464_21_n_936),
       .C (add_464_21_n_915), .Q (add_464_21_n_728));
  ON21X1 add_464_21_g1065(.A (add_464_21_n_874), .B (add_464_21_n_860),
       .C (add_464_21_n_852), .Q (add_464_21_n_729));
  AND2X1 add_464_21_g1066(.A (add_464_21_n_765), .B (add_464_21_n_768),
       .Q (add_464_21_n_730));
  INX1 add_464_21_g1068(.A (add_464_21_n_753), .Q (add_464_21_n_754));
  ON21X1 add_464_21_g1069(.A (add_464_21_n_922), .B (add_464_21_n_931),
       .C (add_464_21_n_912), .Q (add_464_21_n_755));
  ON21X1 add_464_21_g1070(.A (add_464_21_n_938), .B (add_464_21_n_933),
       .C (add_464_21_n_916), .Q (add_464_21_n_756));
  ON21X1 add_464_21_g1071(.A (add_464_21_n_920), .B (add_464_21_n_923),
       .C (add_464_21_n_914), .Q (add_464_21_n_757));
  AND2X1 add_464_21_g1072(.A (add_464_21_n_812), .B (add_464_21_n_939),
       .Q (add_464_21_n_745));
  ON21X1 add_464_21_g1073(.A (add_464_21_n_867), .B (add_464_21_n_872),
       .C (add_464_21_n_853), .Q (add_464_21_n_746));
  NA2X1 add_464_21_g1074(.A (add_464_21_n_769), .B (add_464_21_n_877),
       .Q (add_464_21_n_747));
  AND2X1 add_464_21_g1075(.A (add_464_21_n_807), .B (add_464_21_n_812),
       .Q (add_464_21_n_748));
  AND2X1 add_464_21_g1076(.A (add_464_21_n_811), .B (add_464_21_n_944),
       .Q (add_464_21_n_749));
  ON21X1 add_464_21_g1077(.A (add_464_21_n_918), .B (add_464_21_n_927),
       .C (add_464_21_n_917), .Q (add_464_21_n_750));
  ON21X1 add_464_21_g1078(.A (add_464_21_n_935), .B (add_464_21_n_928),
       .C (add_464_21_n_911), .Q (add_464_21_n_751));
  ON21X1 add_464_21_g1079(.A (add_464_21_n_929), .B (add_464_21_n_921),
       .C (add_464_21_n_913), .Q (add_464_21_n_752));
  NA2X1 add_464_21_g1080(.A (add_464_21_n_808), .B (add_464_21_n_811),
       .Q (add_464_21_n_753));
  NO2I1X1 add_464_21_g1081(.B (add_464_21_n_867), .AN
       (add_464_21_n_853), .Q (add_464_21_n_772));
  NA2X1 add_464_21_g1082(.A (add_464_21_n_865), .B (add_464_21_n_861),
       .Q (add_464_21_n_775));
  NA2I1X1 add_464_21_g1083(.B (add_464_21_n_876), .AN
       (add_464_21_n_864), .Q (add_464_21_n_777));
  NO2I1X1 add_464_21_g1084(.B (add_464_21_n_850), .AN
       (add_464_21_n_871), .Q (add_464_21_n_779));
  AND2X1 add_464_21_g1085(.A (add_464_21_n_868), .B (add_464_21_n_848),
       .Q (add_464_21_n_782));
  NO2I1X1 add_464_21_g1086(.B (add_464_21_n_873), .AN
       (add_464_21_n_851), .Q (add_464_21_n_785));
  AND2X2 add_464_21_g1087(.A (add_464_21_n_871), .B (add_464_21_n_878),
       .Q (add_464_21_n_765));
  NO2X1 add_464_21_g1088(.A (add_464_21_n_873), .B (add_464_21_n_880),
       .Q (add_464_21_n_766));
  NA2X1 add_464_21_g1089(.A (add_464_21_n_881), .B (add_464_21_n_856),
       .Q (add_464_21_n_788));
  NO2I1X1 add_464_21_g1090(.B (add_464_21_n_863), .AN
       (add_464_21_n_878), .Q (add_464_21_n_790));
  NO2I1X1 add_464_21_g1091(.B (add_464_21_n_870), .AN
       (add_464_21_n_860), .Q (add_464_21_n_791));
  AND2X1 add_464_21_g1092(.A (add_464_21_n_879), .B (add_464_21_n_858),
       .Q (add_464_21_n_793));
  NA2I1X1 add_464_21_g1093(.B (add_464_21_n_852), .AN
       (add_464_21_n_874), .Q (add_464_21_n_795));
  NA2X1 add_464_21_g1094(.A (add_464_21_n_877), .B (add_464_21_n_855),
       .Q (add_464_21_n_798));
  NO2I1X1 add_464_21_g1095(.B (add_464_21_n_875), .AN
       (add_464_21_n_949), .Q (add_464_21_n_767));
  NA2I1X1 add_464_21_g1096(.B (add_464_21_n_849), .AN
       (add_464_21_n_866), .Q (add_464_21_n_801));
  NA2I1X1 add_464_21_g1097(.B (add_464_21_n_854), .AN
       (add_464_21_n_875), .Q (add_464_21_n_804));
  NO2X1 add_464_21_g1098(.A (add_464_21_n_870), .B (add_464_21_n_874),
       .Q (add_464_21_n_768));
  NO2X1 add_464_21_g1099(.A (add_464_21_n_943), .B (add_464_21_n_867),
       .Q (add_464_21_n_769));
  NO2X1 add_464_21_g1100(.A (add_464_21_n_864), .B (add_464_21_n_936),
       .Q (add_464_21_n_770));
  NO2X1 add_464_21_g1101(.A (add_464_21_n_882), .B (add_464_21_n_866),
       .Q (add_464_21_n_771));
  AND2X1 add_464_21_g1102(.A (add_464_21_n_948), .B (add_464_21_n_933),
       .Q (add_464_21_n_813));
  NO2I1X1 add_464_21_g1103(.B (add_464_21_n_920), .AN
       (add_464_21_n_914), .Q (add_464_21_n_815));
  NO2I1X1 add_464_21_g1104(.B (add_464_21_n_922), .AN
       (add_464_21_n_912), .Q (add_464_21_n_818));
  NO2X1 add_464_21_g1105(.A (add_464_21_n_922), .B (add_464_21_n_940),
       .Q (add_464_21_n_807));
  NO2X1 add_464_21_g1106(.A (add_464_21_n_920), .B (add_464_21_n_945),
       .Q (add_464_21_n_808));
  AND2X1 add_464_21_g1107(.A (add_464_21_n_944), .B (add_464_21_n_923),
       .Q (add_464_21_n_821));
  AND2X1 add_464_21_g1108(.A (add_464_21_n_939), .B (add_464_21_n_931),
       .Q (add_464_21_n_823));
  AND2X1 add_464_21_g1109(.A (add_464_21_n_946), .B (add_464_21_n_918),
       .Q (add_464_21_n_825));
  AND2X1 add_464_21_g1110(.A (add_464_21_n_941), .B (add_464_21_n_929),
       .Q (add_464_21_n_827));
  NO2I1X1 add_464_21_g1111(.B (add_464_21_n_943), .AN
       (add_464_21_n_872), .Q (add_464_21_n_829));
  AND2X1 add_464_21_g1112(.A (add_464_21_n_949), .B (add_464_21_n_925),
       .Q (add_464_21_n_830));
  NA2I1X1 add_464_21_g1113(.B (add_464_21_n_917), .AN
       (add_464_21_n_927), .Q (add_464_21_n_832));
  NA2I1X1 add_464_21_g1114(.B (add_464_21_n_913), .AN
       (add_464_21_n_921), .Q (add_464_21_n_835));
  NO2I1X1 add_464_21_g1115(.B (add_464_21_n_938), .AN
       (add_464_21_n_916), .Q (add_464_21_n_838));
  NO2I1X1 add_464_21_g1116(.B (add_464_21_n_938), .AN
       (add_464_21_n_948), .Q (add_464_21_n_809));
  NA2I1X1 add_464_21_g1117(.B (add_464_21_n_911), .AN
       (add_464_21_n_935), .Q (add_464_21_n_841));
  NA2I1X1 add_464_21_g1118(.B (add_464_21_n_915), .AN
       (add_464_21_n_936), .Q (add_464_21_n_844));
  NO2I1X1 add_464_21_g1119(.B (add_464_21_n_937), .AN
       (add_464_21_n_928), .Q (add_464_21_n_846));
  NO2X1 add_464_21_g1120(.A (add_464_21_n_937), .B (add_464_21_n_935),
       .Q (add_464_21_n_810));
  NO2X1 add_464_21_g1121(.A (add_464_21_n_942), .B (add_464_21_n_921),
       .Q (add_464_21_n_811));
  NO2X1 add_464_21_g1122(.A (add_464_21_n_947), .B (add_464_21_n_927),
       .Q (add_464_21_n_812));
  INX1 add_464_21_g1123(.A (add_464_21_n_856), .Q (add_464_21_n_857));
  INX1 add_464_21_g1124(.A (add_464_21_n_858), .Q (add_464_21_n_859));
  INX1 add_464_21_g1125(.A (add_464_21_n_861), .Q (add_464_21_n_862));
  INX1 add_464_21_g1126(.A (add_464_21_n_869), .Q (add_464_21_n_868));
  INX1 add_464_21_g1127(.A (add_464_21_n_880), .Q (add_464_21_n_879));
  INX1 add_464_21_g1128(.A (add_464_21_n_882), .Q (add_464_21_n_881));
  NA2X1 add_464_21_g1129(.A (n_7680), .B (program_counter[3]), .Q
       (add_464_21_n_848));
  NA2X1 add_464_21_g1130(.A (n_7689), .B (program_counter[13]), .Q
       (add_464_21_n_849));
  AND2X1 add_464_21_g1131(.A (n_7683), .B (program_counter[19]), .Q
       (add_464_21_n_850));
  NA2X1 add_464_21_g1132(.A (n_7687), .B (program_counter[15]), .Q
       (add_464_21_n_851));
  NA2X1 add_464_21_g1133(.A (n_7685), .B (program_counter[17]), .Q
       (add_464_21_n_852));
  NA2X1 add_464_21_g1134(.A (n_7672), .B (program_counter[29]), .Q
       (add_464_21_n_853));
  NA2X1 add_464_21_g1135(.A (n_7691), .B (program_counter[11]), .Q
       (add_464_21_n_854));
  NA2X1 add_464_21_g1136(.A (n_7671), .B (program_counter[30]), .Q
       (add_464_21_n_855));
  NA2X1 add_464_21_g1137(.A (n_7690), .B (program_counter[12]), .Q
       (add_464_21_n_856));
  NA2X1 add_464_21_g1138(.A (n_7688), .B (program_counter[14]), .Q
       (add_464_21_n_858));
  NA2X1 add_464_21_g1139(.A (n_7686), .B (program_counter[16]), .Q
       (add_464_21_n_860));
  NA2X1 add_464_21_g1140(.A (n_7681), .B (program_counter[2]), .Q
       (add_464_21_n_861));
  AND2X1 add_464_21_g1141(.A (n_7684), .B (program_counter[18]), .Q
       (add_464_21_n_863));
  NO2X1 add_464_21_g1142(.A (n_2437), .B (program_counter[4]), .Q
       (add_464_21_n_864));
  OR2X1 add_464_21_g1143(.A (n_7681), .B (program_counter[2]), .Q
       (add_464_21_n_865));
  NO2X1 add_464_21_g1144(.A (n_7689), .B (program_counter[13]), .Q
       (add_464_21_n_866));
  NO2X1 add_464_21_g1145(.A (n_7672), .B (program_counter[29]), .Q
       (add_464_21_n_867));
  NO2X1 add_464_21_g1146(.A (n_7680), .B (program_counter[3]), .Q
       (add_464_21_n_869));
  NO2X1 add_464_21_g1147(.A (n_7686), .B (program_counter[16]), .Q
       (add_464_21_n_870));
  OR2X2 add_464_21_g1148(.A (n_7683), .B (program_counter[19]), .Q
       (add_464_21_n_871));
  NA2X1 add_464_21_g1149(.A (n_7673), .B (program_counter[28]), .Q
       (add_464_21_n_872));
  NO2X1 add_464_21_g1150(.A (n_7687), .B (program_counter[15]), .Q
       (add_464_21_n_873));
  NO2X1 add_464_21_g1151(.A (n_7685), .B (program_counter[17]), .Q
       (add_464_21_n_874));
  NO2X1 add_464_21_g1152(.A (n_7691), .B (program_counter[11]), .Q
       (add_464_21_n_875));
  NA2X1 add_464_21_g1153(.A (n_2437), .B (program_counter[4]), .Q
       (add_464_21_n_876));
  OR2X1 add_464_21_g1154(.A (n_7671), .B (program_counter[30]), .Q
       (add_464_21_n_877));
  OR2X2 add_464_21_g1155(.A (n_7684), .B (program_counter[18]), .Q
       (add_464_21_n_878));
  NO2X1 add_464_21_g1156(.A (n_7688), .B (program_counter[14]), .Q
       (add_464_21_n_880));
  NO2X1 add_464_21_g1157(.A (n_7690), .B (program_counter[12]), .Q
       (add_464_21_n_882));
  INX1 add_464_21_g1158(.A (add_464_21_n_918), .Q (add_464_21_n_919));
  INX1 add_464_21_g1159(.A (add_464_21_n_923), .Q (add_464_21_n_924));
  INX1 add_464_21_g1160(.A (add_464_21_n_925), .Q (add_464_21_n_926));
  INX1 add_464_21_g1161(.A (add_464_21_n_929), .Q (add_464_21_n_930));
  INX1 add_464_21_g1162(.A (add_464_21_n_931), .Q (add_464_21_n_932));
  INX1 add_464_21_g1163(.A (add_464_21_n_933), .Q (add_464_21_n_934));
  INX1 add_464_21_g1164(.A (add_464_21_n_940), .Q (add_464_21_n_939));
  INX1 add_464_21_g1165(.A (add_464_21_n_942), .Q (add_464_21_n_941));
  INX1 add_464_21_g1166(.A (add_464_21_n_945), .Q (add_464_21_n_944));
  INX1 add_464_21_g1167(.A (add_464_21_n_947), .Q (add_464_21_n_946));
  NA2X1 add_464_21_g1168(.A (n_8261), .B (program_counter[9]), .Q
       (add_464_21_n_911));
  NA2X1 add_464_21_g1169(.A (n_7678), .B (program_counter[23]), .Q
       (add_464_21_n_912));
  NA2X1 add_464_21_g1170(.A (n_7676), .B (program_counter[25]), .Q
       (add_464_21_n_913));
  NA2X1 add_464_21_g1171(.A (n_7674), .B (program_counter[27]), .Q
       (add_464_21_n_914));
  NA2X1 add_464_21_g1172(.A (n_8257), .B (program_counter[5]), .Q
       (add_464_21_n_915));
  NA2X1 add_464_21_g1173(.A (n_8259), .B (program_counter[7]), .Q
       (add_464_21_n_916));
  NA2X1 add_464_21_g1174(.A (n_7693), .B (program_counter[21]), .Q
       (add_464_21_n_917));
  NA2X1 add_464_21_g1175(.A (n_7670), .B (program_counter[20]), .Q
       (add_464_21_n_918));
  NO2X1 add_464_21_g1176(.A (n_7674), .B (program_counter[27]), .Q
       (add_464_21_n_920));
  NO2X1 add_464_21_g1177(.A (n_7676), .B (program_counter[25]), .Q
       (add_464_21_n_921));
  NO2X1 add_464_21_g1178(.A (n_7678), .B (program_counter[23]), .Q
       (add_464_21_n_922));
  NA2X1 add_464_21_g1179(.A (n_7675), .B (program_counter[26]), .Q
       (add_464_21_n_923));
  NA2X1 add_464_21_g1180(.A (n_8262), .B (program_counter[10]), .Q
       (add_464_21_n_925));
  NO2X1 add_464_21_g1181(.A (n_7693), .B (program_counter[21]), .Q
       (add_464_21_n_927));
  NA2X1 add_464_21_g1182(.A (n_8260), .B (program_counter[8]), .Q
       (add_464_21_n_928));
  NA2X1 add_464_21_g1183(.A (n_7677), .B (program_counter[24]), .Q
       (add_464_21_n_929));
  NA2X1 add_464_21_g1184(.A (n_7669), .B (program_counter[22]), .Q
       (add_464_21_n_931));
  NA2X1 add_464_21_g1185(.A (n_8258), .B (program_counter[6]), .Q
       (add_464_21_n_933));
  NO2X1 add_464_21_g1186(.A (n_8261), .B (program_counter[9]), .Q
       (add_464_21_n_935));
  NO2X1 add_464_21_g1187(.A (n_8257), .B (program_counter[5]), .Q
       (add_464_21_n_936));
  NO2X1 add_464_21_g1188(.A (n_8260), .B (program_counter[8]), .Q
       (add_464_21_n_937));
  NO2X1 add_464_21_g1189(.A (n_8259), .B (program_counter[7]), .Q
       (add_464_21_n_938));
  NO2X1 add_464_21_g1190(.A (n_7669), .B (program_counter[22]), .Q
       (add_464_21_n_940));
  NO2X1 add_464_21_g1191(.A (n_7677), .B (program_counter[24]), .Q
       (add_464_21_n_942));
  NO2X1 add_464_21_g1192(.A (n_7673), .B (program_counter[28]), .Q
       (add_464_21_n_943));
  NO2X1 add_464_21_g1193(.A (n_7675), .B (program_counter[26]), .Q
       (add_464_21_n_945));
  NO2X1 add_464_21_g1194(.A (n_7670), .B (program_counter[20]), .Q
       (add_464_21_n_947));
  OR2X1 add_464_21_g1195(.A (n_8258), .B (program_counter[6]), .Q
       (add_464_21_n_948));
  OR2X1 add_464_21_g1196(.A (n_8262), .B (program_counter[10]), .Q
       (add_464_21_n_949));
  AND2X1 add_464_21_g1198(.A (add_464_21_n_767), .B (add_464_21_n_810),
       .Q (add_464_21_n_731));
  EN3X1 add_464_21_g1200(.A (add_464_21_n_602), .B (n_8263), .C
       (program_counter[31]), .Q (n_7765));
  AO321X1 add_464_21_g1202(.A (add_464_21_n_881), .B
       (add_464_21_n_731), .C (add_464_21_n_653), .D
       (add_464_21_n_881), .E (add_464_21_n_702), .F
       (add_464_21_n_857), .Q (add_464_21_n_639));
  AO321X1 add_464_21_g1204(.A (add_464_21_n_949), .B
       (add_464_21_n_810), .C (add_464_21_n_653), .D
       (add_464_21_n_949), .E (add_464_21_n_751), .F
       (add_464_21_n_926), .Q (add_464_21_n_643));
  AND2X1 add_464_21_g1206(.A (add_464_21_n_730), .B (add_464_21_n_748),
       .Q (add_464_21_n_708));
  MU2IX1 inc_ADD_UNS_OP_5_g3281(.S (inc_ADD_UNS_OP_5_n_3387), .IN0
       (n_7376), .IN1 (inc_ADD_UNS_OP_5_n_3752), .Q (n_7435));
  NO2X4 inc_ADD_UNS_OP_5_g3283(.A (inc_ADD_UNS_OP_5_n_3387), .B
       (inc_ADD_UNS_OP_5_n_3752), .Q (inc_ADD_UNS_OP_5_n_3370));
  NA2X2 inc_ADD_UNS_OP_5_g3291(.A (inc_ADD_UNS_OP_5_n_3411), .B
       (n_7377), .Q (inc_ADD_UNS_OP_5_n_3387));
  NO2X2 inc_ADD_UNS_OP_5_g3294(.A (inc_ADD_UNS_OP_5_n_3415), .B
       (inc_ADD_UNS_OP_5_n_3792), .Q (inc_ADD_UNS_OP_5_n_3392));
  MU2IX1 inc_ADD_UNS_OP_5_g3297(.S (inc_ADD_UNS_OP_5_n_3424), .IN0
       (csr_minstret[53]), .IN1 (inc_ADD_UNS_OP_5_n_3832), .Q (n_7412));
  NO2X4 inc_ADD_UNS_OP_5_g3299(.A (inc_ADD_UNS_OP_5_n_3424), .B
       (inc_ADD_UNS_OP_5_n_3832), .Q (inc_ADD_UNS_OP_5_n_3400));
  MU2IX1 inc_ADD_UNS_OP_5_g3302(.S (inc_ADD_UNS_OP_5_n_3430), .IN0
       (n_7378), .IN1 (inc_ADD_UNS_OP_5_n_3742), .Q (n_7437));
  NO2X4 inc_ADD_UNS_OP_5_g3304(.A (inc_ADD_UNS_OP_5_n_3430), .B
       (inc_ADD_UNS_OP_5_n_3742), .Q (inc_ADD_UNS_OP_5_n_3411));
  NA2X4 inc_ADD_UNS_OP_5_g3305(.A (inc_ADD_UNS_OP_5_n_3438), .B
       (csr_minstret[61]), .Q (inc_ADD_UNS_OP_5_n_3415));
  MU2IX1 inc_ADD_UNS_OP_5_g3306(.S (inc_ADD_UNS_OP_5_n_3432), .IN0
       (csr_minstret[32]), .IN1 (inc_ADD_UNS_OP_5_n_3834), .Q (n_7433));
  NO2X4 inc_ADD_UNS_OP_5_g3309(.A (inc_ADD_UNS_OP_5_n_3432), .B
       (inc_ADD_UNS_OP_5_n_3834), .Q (inc_ADD_UNS_OP_5_n_3421));
  NA2X4 inc_ADD_UNS_OP_5_g3310(.A (inc_ADD_UNS_OP_5_n_3447), .B
       (csr_minstret[52]), .Q (inc_ADD_UNS_OP_5_n_3424));
  NA2X4 inc_ADD_UNS_OP_5_g3314(.A (inc_ADD_UNS_OP_5_n_3453), .B
       (n_7379), .Q (inc_ADD_UNS_OP_5_n_3430));
  NA2X4 inc_ADD_UNS_OP_5_g3315(.A (inc_ADD_UNS_OP_5_n_3435), .B
       (inc_ADD_UNS_OP_5_n_3711), .Q (inc_ADD_UNS_OP_5_n_3432));
  BUX1 inc_ADD_UNS_OP_5_g3317(.A (inc_ADD_UNS_OP_5_n_3453), .Q
       (inc_ADD_UNS_OP_5_n_3435));
  NO2X4 inc_ADD_UNS_OP_5_g3319(.A (inc_ADD_UNS_OP_5_n_3445), .B
       (inc_ADD_UNS_OP_5_n_3785), .Q (inc_ADD_UNS_OP_5_n_3438));
  MU2IX1 inc_ADD_UNS_OP_5_g3321(.S (inc_ADD_UNS_OP_5_n_3463), .IN0
       (csr_minstret[51]), .IN1 (inc_ADD_UNS_OP_5_n_3824), .Q (n_7414));
  NO2X4 inc_ADD_UNS_OP_5_g3325(.A (inc_ADD_UNS_OP_5_n_3463), .B
       (inc_ADD_UNS_OP_5_n_3824), .Q (inc_ADD_UNS_OP_5_n_3447));
  MU2IX1 inc_ADD_UNS_OP_5_g3326(.S (inc_ADD_UNS_OP_5_n_3470), .IN0
       (n_7380), .IN1 (inc_ADD_UNS_OP_5_n_3775), .Q (n_7439));
  NO2X4 inc_ADD_UNS_OP_5_g3328(.A (inc_ADD_UNS_OP_5_n_3470), .B
       (inc_ADD_UNS_OP_5_n_3775), .Q (inc_ADD_UNS_OP_5_n_3453));
  NA2X4 inc_ADD_UNS_OP_5_g3329(.A (inc_ADD_UNS_OP_5_n_3476), .B
       (csr_minstret[59]), .Q (inc_ADD_UNS_OP_5_n_3445));
  NA2X4 inc_ADD_UNS_OP_5_g3333(.A (inc_ADD_UNS_OP_5_n_3482), .B
       (csr_minstret[50]), .Q (inc_ADD_UNS_OP_5_n_3463));
  MU2IX1 inc_ADD_UNS_OP_5_g3336(.S (inc_ADD_UNS_OP_5_n_3494), .IN0
       (csr_minstret[58]), .IN1 (inc_ADD_UNS_OP_5_n_3803), .Q (n_7407));
  NA2X1 inc_ADD_UNS_OP_5_g3337(.A (inc_ADD_UNS_OP_5_n_3474), .B
       (inc_ADD_UNS_OP_5_n_3695), .Q (inc_ADD_UNS_OP_5_n_3469));
  NA2X4 inc_ADD_UNS_OP_5_g3338(.A (inc_ADD_UNS_OP_5_n_3490), .B
       (n_7381), .Q (inc_ADD_UNS_OP_5_n_3470));
  NO2X4 inc_ADD_UNS_OP_5_g3342(.A (inc_ADD_UNS_OP_5_n_3494), .B
       (inc_ADD_UNS_OP_5_n_3803), .Q (inc_ADD_UNS_OP_5_n_3476));
  MU2IX1 inc_ADD_UNS_OP_5_g3343(.S (inc_ADD_UNS_OP_5_n_3499), .IN0
       (csr_minstret[49]), .IN1 (inc_ADD_UNS_OP_5_n_3826), .Q (n_7416));
  NO2X4 inc_ADD_UNS_OP_5_g3345(.A (inc_ADD_UNS_OP_5_n_3499), .B
       (inc_ADD_UNS_OP_5_n_3826), .Q (inc_ADD_UNS_OP_5_n_3482));
  MU2IX1 inc_ADD_UNS_OP_5_g3346(.S (inc_ADD_UNS_OP_5_n_3505), .IN0
       (n_8571), .IN1 (inc_ADD_UNS_OP_5_n_3756), .Q (n_7441));
  BUX1 inc_ADD_UNS_OP_5_g3348(.A (inc_ADD_UNS_OP_5_n_3490), .Q
       (inc_ADD_UNS_OP_5_n_3474));
  NO2X4 inc_ADD_UNS_OP_5_g3349(.A (inc_ADD_UNS_OP_5_n_3505), .B
       (inc_ADD_UNS_OP_5_n_3756), .Q (inc_ADD_UNS_OP_5_n_3490));
  NA2X4 inc_ADD_UNS_OP_5_g3350(.A (inc_ADD_UNS_OP_5_n_3509), .B
       (csr_minstret[57]), .Q (inc_ADD_UNS_OP_5_n_3494));
  NA2X4 inc_ADD_UNS_OP_5_g3353(.A (inc_ADD_UNS_OP_5_n_3515), .B
       (csr_minstret[48]), .Q (inc_ADD_UNS_OP_5_n_3499));
  MU2IX1 inc_ADD_UNS_OP_5_g3356(.S (inc_ADD_UNS_OP_5_n_3527), .IN0
       (csr_minstret[56]), .IN1 (inc_ADD_UNS_OP_5_n_3795), .Q (n_7409));
  NA2X4 inc_ADD_UNS_OP_5_g3357(.A (inc_ADD_UNS_OP_5_n_3522), .B
       (n_7383), .Q (inc_ADD_UNS_OP_5_n_3505));
  NO2X2 inc_ADD_UNS_OP_5_g3360(.A (inc_ADD_UNS_OP_5_n_3527), .B
       (inc_ADD_UNS_OP_5_n_3795), .Q (inc_ADD_UNS_OP_5_n_3509));
  MU2IX1 inc_ADD_UNS_OP_5_g3361(.S (inc_ADD_UNS_OP_5_n_3531), .IN0
       (csr_minstret[47]), .IN1 (inc_ADD_UNS_OP_5_n_3838), .Q (n_7418));
  NO2X4 inc_ADD_UNS_OP_5_g3363(.A (inc_ADD_UNS_OP_5_n_3531), .B
       (inc_ADD_UNS_OP_5_n_3838), .Q (inc_ADD_UNS_OP_5_n_3515));
  MU2IX1 inc_ADD_UNS_OP_5_g3364(.S (inc_ADD_UNS_OP_5_n_3538), .IN0
       (n_7384), .IN1 (inc_ADD_UNS_OP_5_n_3746), .Q (n_7443));
  MU2IX1 inc_ADD_UNS_OP_5_g3365(.S (inc_ADD_UNS_OP_5_n_3530), .IN0
       (csr_minstret[55]), .IN1 (inc_ADD_UNS_OP5492_3_n_2608), .Q
       (n_7410));
  NO2X4 inc_ADD_UNS_OP_5_g3367(.A (inc_ADD_UNS_OP_5_n_3538), .B
       (inc_ADD_UNS_OP_5_n_3746), .Q (inc_ADD_UNS_OP_5_n_3522));
  OR6X2 inc_ADD_UNS_OP_5_g3368(.A (inc_ADD_UNS_OP_5_n_3574), .B
       (inc_ADD_UNS_OP_5_n_3703), .C (inc_ADD_UNS_OP_5_n_3800), .D
       (inc_ADD_UNS_OP_5_n_3791), .E (inc_ADD_UNS_OP5492_3_n_2613), .F
       (inc_ADD_UNS_OP5492_3_n_2608), .Q (inc_ADD_UNS_OP_5_n_3527));
  NA2X1 inc_ADD_UNS_OP_5_g3370(.A (inc_ADD_UNS_OP_5_n_3536), .B
       (inc_ADD_UNS_OP_5_n_3704), .Q (inc_ADD_UNS_OP_5_n_3530));
  NA2X4 inc_ADD_UNS_OP_5_g3371(.A (inc_ADD_UNS_OP_5_n_3536), .B
       (csr_minstret[46]), .Q (inc_ADD_UNS_OP_5_n_3531));
  NA2X4 inc_ADD_UNS_OP_5_g3375(.A (inc_ADD_UNS_OP_5_n_3541), .B
       (n_7385), .Q (inc_ADD_UNS_OP_5_n_3538));
  MU2IX1 inc_ADD_UNS_OP_5_g3377(.S (inc_ADD_UNS_OP_5_n_3556), .IN0
       (csr_minstret[45]), .IN1 (inc_ADD_UNS_OP5492_3_n_2613), .Q
       (n_7420));
  AND6X2 inc_ADD_UNS_OP_5_g3379(.A (inc_ADD_UNS_OP_5_n_3611), .B
       (csr_minstret[41]), .C (csr_minstret[43]), .D
       (csr_minstret[42]), .E (csr_minstret[44]), .F
       (csr_minstret[45]), .Q (inc_ADD_UNS_OP_5_n_3536));
  MU2IX1 inc_ADD_UNS_OP_5_g3380(.S (inc_ADD_UNS_OP_5_n_3559), .IN0
       (n_7386), .IN1 (inc_ADD_UNS_OP_5_n_3760), .Q (n_7445));
  NO2X4 inc_ADD_UNS_OP_5_g3381(.A (inc_ADD_UNS_OP_5_n_3559), .B
       (inc_ADD_UNS_OP_5_n_3760), .Q (inc_ADD_UNS_OP_5_n_3541));
  MU2IX1 inc_ADD_UNS_OP_5_g3382(.S (inc_ADD_UNS_OP_5_n_3567), .IN0
       (csr_minstret[44]), .IN1 (inc_ADD_UNS_OP_5_n_3791), .Q (n_7421));
  NA3X1 inc_ADD_UNS_OP_5_g3383(.A (inc_ADD_UNS_OP_5_n_3573), .B
       (csr_minstret[43]), .C (csr_minstret[44]), .Q
       (inc_ADD_UNS_OP_5_n_3556));
  NA2X4 inc_ADD_UNS_OP_5_g3385(.A (inc_ADD_UNS_OP_5_n_3581), .B
       (n_7387), .Q (inc_ADD_UNS_OP_5_n_3559));
  MU2IX1 inc_ADD_UNS_OP_5_g3388(.S (inc_ADD_UNS_OP_5_n_3574), .IN0
       (csr_minstret[43]), .IN1 (inc_ADD_UNS_OP_5_n_3800), .Q (n_7422));
  NA2X1 inc_ADD_UNS_OP_5_g3389(.A (inc_ADD_UNS_OP_5_n_3573), .B
       (csr_minstret[43]), .Q (inc_ADD_UNS_OP_5_n_3567));
  MU2IX1 inc_ADD_UNS_OP_5_g3392(.S (inc_ADD_UNS_OP_5_n_3583), .IN0
       (n_7388), .IN1 (inc_ADD_UNS_OP_5_n_3748), .Q (n_7447));
  INX1 inc_ADD_UNS_OP_5_g3393(.A (inc_ADD_UNS_OP_5_n_3574), .Q
       (inc_ADD_UNS_OP_5_n_3573));
  BUX1 inc_ADD_UNS_OP_5_g3398(.A (inc_ADD_UNS_OP_5_n_3581), .Q
       (inc_ADD_UNS_OP_5_n_3580));
  NO2X4 inc_ADD_UNS_OP_5_g3399(.A (inc_ADD_UNS_OP_5_n_3590), .B
       (inc_ADD_UNS_OP_5_n_3748), .Q (inc_ADD_UNS_OP_5_n_3581));
  BUX1 inc_ADD_UNS_OP_5_g3400(.A (inc_ADD_UNS_OP_5_n_3590), .Q
       (inc_ADD_UNS_OP_5_n_3583));
  MU2IX1 inc_ADD_UNS_OP_5_g3401(.S (inc_ADD_UNS_OP_5_n_3597), .IN0
       (csr_minstret[42]), .IN1 (inc_ADD_UNS_OP_5_n_3808), .Q (n_7423));
  OR6X2 inc_ADD_UNS_OP_5_g3402(.A (inc_ADD_UNS_OP_5_n_3637), .B
       (inc_ADD_UNS_OP_5_n_3798), .C (inc_ADD_UNS_OP_5_n_3815), .D
       (inc_ADD_UNS_OP_5_n_3789), .E (inc_ADD_UNS_OP_5_n_3812), .F
       (inc_ADD_UNS_OP_5_n_3808), .Q (inc_ADD_UNS_OP_5_n_3574));
  NA2X4 inc_ADD_UNS_OP_5_g3404(.A (inc_ADD_UNS_OP_5_n_3606), .B
       (n_7389), .Q (inc_ADD_UNS_OP_5_n_3590));
  MU2IX1 inc_ADD_UNS_OP_5_g3408(.S (inc_ADD_UNS_OP_5_n_3616), .IN0
       (n_8622), .IN1 (inc_ADD_UNS_OP_5_n_3768), .Q (n_7449));
  BUX1 inc_ADD_UNS_OP_5_g3410(.A (inc_ADD_UNS_OP_5_n_3606), .Q
       (inc_ADD_UNS_OP_5_n_3605));
  NO2X4 inc_ADD_UNS_OP_5_g3411(.A (inc_ADD_UNS_OP_5_n_3616), .B
       (inc_ADD_UNS_OP_5_n_3768), .Q (inc_ADD_UNS_OP_5_n_3606));
  EN2X1 inc_ADD_UNS_OP_5_g3412(.A (inc_ADD_UNS_OP_5_n_3614), .B
       (inc_ADD_UNS_OP_5_n_3815), .Q (n_7425));
  AND6X2 inc_ADD_UNS_OP_5_g3413(.A (inc_ADD_UNS_OP_5_n_3651), .B
       (csr_minstret[36]), .C (csr_minstret[38]), .D
       (csr_minstret[37]), .E (csr_minstret[39]), .F
       (csr_minstret[40]), .Q (inc_ADD_UNS_OP_5_n_3611));
  HAX1 inc_ADD_UNS_OP_5_g3415(.A (inc_ADD_UNS_OP_5_n_3628), .B
       (csr_minstret[39]), .S (n_7426), .CO (inc_ADD_UNS_OP_5_n_3614));
  NA2X4 inc_ADD_UNS_OP_5_g3416(.A (inc_ADD_UNS_OP_5_n_3622), .B
       (n_7391), .Q (inc_ADD_UNS_OP_5_n_3616));
  MU2IX1 inc_ADD_UNS_OP_5_g3418(.S (inc_ADD_UNS_OP_5_n_3631), .IN0
       (n_7392), .IN1 (inc_ADD_UNS_OP_5_n_3766), .Q (n_7451));
  BUX1 inc_ADD_UNS_OP_5_g3419(.A (inc_ADD_UNS_OP_5_n_3622), .Q
       (inc_ADD_UNS_OP_5_n_3621));
  NO2X4 inc_ADD_UNS_OP_5_g3420(.A (inc_ADD_UNS_OP_5_n_3631), .B
       (inc_ADD_UNS_OP_5_n_3766), .Q (inc_ADD_UNS_OP_5_n_3622));
  EN2X1 inc_ADD_UNS_OP_5_g3421(.A (inc_ADD_UNS_OP_5_n_3637), .B
       (csr_minstret[38]), .Q (n_7427));
  NO2X1 inc_ADD_UNS_OP_5_g3422(.A (inc_ADD_UNS_OP_5_n_3637), .B
       (inc_ADD_UNS_OP_5_n_3798), .Q (inc_ADD_UNS_OP_5_n_3628));
  NA2X4 inc_ADD_UNS_OP_5_g3424(.A (inc_ADD_UNS_OP_5_n_3643), .B
       (n_7393), .Q (inc_ADD_UNS_OP_5_n_3631));
  EO2X1 inc_ADD_UNS_OP_5_g3426(.A (inc_ADD_UNS_OP_5_n_3641), .B
       (csr_minstret[37]), .Q (n_7428));
  NA6X4 inc_ADD_UNS_OP_5_g3427(.A (inc_ADD_UNS_OP_5_n_3665), .B
       (inc_ADD_UNS_OP_5_n_3686), .C (n_7397), .D (n_8354), .E
       (csr_minstret[36]), .F (csr_minstret[37]), .Q
       (inc_ADD_UNS_OP_5_n_3637));
  MU2IX1 inc_ADD_UNS_OP_5_g3428(.S (inc_ADD_UNS_OP_5_n_3645), .IN0
       (inc_ADD_UNS_OP_5_n_3750), .IN1 (n_7394), .Q (n_7453));
  HAX1 inc_ADD_UNS_OP_5_g3429(.A (inc_ADD_UNS_OP_5_n_3651), .B
       (csr_minstret[36]), .S (n_7429), .CO (inc_ADD_UNS_OP_5_n_3641));
  NO2X4 inc_ADD_UNS_OP_5_g3430(.A (inc_ADD_UNS_OP_5_n_3648), .B
       (inc_ADD_UNS_OP_5_n_3750), .Q (inc_ADD_UNS_OP_5_n_3643));
  INX1 inc_ADD_UNS_OP_5_g3431(.A (inc_ADD_UNS_OP_5_n_3648), .Q
       (inc_ADD_UNS_OP_5_n_3645));
  NA2X4 inc_ADD_UNS_OP_5_g3433(.A (inc_ADD_UNS_OP_5_n_3658), .B
       (n_7395), .Q (inc_ADD_UNS_OP_5_n_3648));
  AND6X2 inc_ADD_UNS_OP_5_g3434(.A (inc_ADD_UNS_OP_5_n_3670), .B
       (inc_ADD_UNS_OP_5_n_3686), .C (n_6238), .D (n_8354), .E
       (n_7398), .F (n_7397), .Q (inc_ADD_UNS_OP_5_n_3651));
  BUX1 inc_ADD_UNS_OP_5_g3435(.A (inc_ADD_UNS_OP_5_n_3658), .Q
       (inc_ADD_UNS_OP_5_n_3655));
  EN2X1 inc_ADD_UNS_OP_5_g3436(.A (inc_ADD_UNS_OP_5_n_3663), .B
       (n_8354), .Q (n_7455));
  AND6X2 inc_ADD_UNS_OP_5_g3437(.A (inc_ADD_UNS_OP_5_n_3676), .B
       (n_6237), .C (n_6238), .D (n_8354), .E (n_7398), .F (n_7397), .Q
       (inc_ADD_UNS_OP_5_n_3658));
  EO2X1 inc_ADD_UNS_OP_5_g3438(.A (inc_ADD_UNS_OP_5_n_3664), .B
       (n_7397), .Q (n_7456));
  NA2X1 inc_ADD_UNS_OP_5_g3439(.A (inc_ADD_UNS_OP_5_n_3664), .B
       (n_7397), .Q (inc_ADD_UNS_OP_5_n_3663));
  BUX1 inc_ADD_UNS_OP_5_g3440(.A (inc_ADD_UNS_OP_5_n_3665), .Q
       (inc_ADD_UNS_OP_5_n_3664));
  HAX2 inc_ADD_UNS_OP_5_g3441(.A (inc_ADD_UNS_OP_5_n_3668), .B
       (n_7398), .S (n_7457), .CO (inc_ADD_UNS_OP_5_n_3665));
  HAX2 inc_ADD_UNS_OP_5_g3442(.A (inc_ADD_UNS_OP_5_n_3670), .B
       (n_6238), .S (n_7458), .CO (inc_ADD_UNS_OP_5_n_3668));
  HAX2 inc_ADD_UNS_OP_5_g3443(.A (inc_ADD_UNS_OP_5_n_3676), .B
       (n_6237), .S (n_7459), .CO (inc_ADD_UNS_OP_5_n_3670));
  NO2I1X4 inc_ADD_UNS_OP_5_g3445(.B (inc_ADD_UNS_OP_5_n_3681), .AN
       (n_6232), .Q (inc_ADD_UNS_OP_5_n_3676));
  EO2X1 inc_ADD_UNS_OP_5_g3447(.A (inc_ADD_UNS_OP_5_n_3684), .B
       (n_7632), .Q (n_7461));
  NA2X4 inc_ADD_UNS_OP_5_g3448(.A (inc_ADD_UNS_OP_5_n_3684), .B
       (n_7632), .Q (inc_ADD_UNS_OP_5_n_3681));
  HAX4 inc_ADD_UNS_OP_5_g3449(.A (inc_ADD_UNS_OP_5_n_3692), .B
       (n_6234), .S (n_7462), .CO (inc_ADD_UNS_OP_5_n_3684));
  AND5X2 inc_ADD_UNS_OP_5_g3450(.A (inc_ADD_UNS_OP_5_n_3697), .B
       (inc_ADD_UNS_OP_5_n_3711), .C (inc_ADD_UNS_OP_5_n_3724), .D
       (inc_ADD_UNS_OP_5_n_3714), .E (inc_ADD_UNS_OP_5_n_3717), .Q
       (inc_ADD_UNS_OP_5_n_3686));
  EN2X0 inc_ADD_UNS_OP_5_g3451(.A (inc_ADD_UNS_OP_5_n_3701), .B
       (n_7633), .Q (n_7463));
  NO2X2 inc_ADD_UNS_OP_5_g3453(.A (inc_ADD_UNS_OP_5_n_3701), .B
       (inc_ADD_UNS_OP_5_n_3733), .Q (inc_ADD_UNS_OP_5_n_3692));
  EO2X1 inc_ADD_UNS_OP_5_g3454(.A (inc_ADD_UNS_OP_5_n_3708), .B
       (n_6235), .Q (n_7464));
  AND2X1 inc_ADD_UNS_OP_5_g3455(.A (inc_ADD_UNS_OP_5_n_3711), .B
       (inc_ADD_UNS_OP_5_n_3714), .Q (inc_ADD_UNS_OP_5_n_3695));
  AND6X2 inc_ADD_UNS_OP_5_g3456(.A (inc_ADD_UNS_OP_5_n_3726), .B
       (n_7384), .C (n_7386), .D (n_7385), .E (n_8571), .F (n_7387), .Q
       (inc_ADD_UNS_OP_5_n_3697));
  NA3X2 inc_ADD_UNS_OP_5_g3457(.A (n_7636), .B (n_6235), .C (n_7883),
       .Q (inc_ADD_UNS_OP_5_n_3701));
  INX1 inc_ADD_UNS_OP_5_g3458(.A (inc_ADD_UNS_OP_5_n_3704), .Q
       (inc_ADD_UNS_OP_5_n_3703));
  AND5X1 inc_ADD_UNS_OP_5_g3459(.A (inc_ADD_UNS_OP_5_n_3721), .B
       (csr_minstret[46]), .C (csr_minstret[47]), .D
       (csr_minstret[53]), .E (csr_minstret[52]), .Q
       (inc_ADD_UNS_OP_5_n_3704));
  HAX1 inc_ADD_UNS_OP_5_g3460(.A (n_7636), .B (n_7883), .S (n_7465),
       .CO (inc_ADD_UNS_OP_5_n_3708));
  AND5X2 inc_ADD_UNS_OP_5_g3461(.A (n_7379), .B (n_7635), .C (n_7376),
       .D (n_7378), .E (n_7377), .Q (inc_ADD_UNS_OP_5_n_3711));
  AND4X1 inc_ADD_UNS_OP_5_g3462(.A (n_7380), .B (n_7381), .C
       (csr_minstret[32]), .D (csr_minstret[33]), .Q
       (inc_ADD_UNS_OP_5_n_3714));
  AND5X1 inc_ADD_UNS_OP_5_g3463(.A (n_7394), .B (n_7395), .C (n_8622),
       .D (n_7389), .E (csr_minstret[35]), .Q
       (inc_ADD_UNS_OP_5_n_3717));
  AND5X1 inc_ADD_UNS_OP_5_g3464(.A (csr_minstret[48]), .B
       (csr_minstret[54]), .C (csr_minstret[50]), .D
       (csr_minstret[49]), .E (csr_minstret[51]), .Q
       (inc_ADD_UNS_OP_5_n_3721));
  AND3X1 inc_ADD_UNS_OP_5_g3465(.A (n_7392), .B (n_7391), .C (n_7393),
       .Q (inc_ADD_UNS_OP_5_n_3724));
  AND3X1 inc_ADD_UNS_OP_5_g3466(.A (n_7383), .B (n_7388), .C
       (csr_minstret[34]), .Q (inc_ADD_UNS_OP_5_n_3726));
  INX1 inc_ADD_UNS_OP_5_g3467(.A (n_7633), .Q
       (inc_ADD_UNS_OP_5_n_3733));
  INX1 inc_ADD_UNS_OP_5_g3468(.A (n_7635), .Q
       (inc_ADD_UNS_OP_5_n_3735));
  INX1 inc_ADD_UNS_OP_5_g3469(.A (n_7378), .Q
       (inc_ADD_UNS_OP_5_n_3742));
  INX1 inc_ADD_UNS_OP_5_g3471(.A (n_7384), .Q
       (inc_ADD_UNS_OP_5_n_3746));
  INX1 inc_ADD_UNS_OP_5_g3472(.A (n_7388), .Q
       (inc_ADD_UNS_OP_5_n_3748));
  INX1 inc_ADD_UNS_OP_5_g3473(.A (n_7394), .Q
       (inc_ADD_UNS_OP_5_n_3750));
  INX1 inc_ADD_UNS_OP_5_g3474(.A (n_7376), .Q
       (inc_ADD_UNS_OP_5_n_3752));
  INX1 inc_ADD_UNS_OP_5_g3476(.A (n_8571), .Q
       (inc_ADD_UNS_OP_5_n_3756));
  INX1 inc_ADD_UNS_OP_5_g3478(.A (n_7386), .Q
       (inc_ADD_UNS_OP_5_n_3760));
  INX1 inc_ADD_UNS_OP_5_g3482(.A (n_8622), .Q
       (inc_ADD_UNS_OP_5_n_3768));
  INX1 inc_ADD_UNS_OP_5_g3485(.A (n_7380), .Q
       (inc_ADD_UNS_OP_5_n_3775));
  INX1 inc_ADD_UNS_OP_5_g3489(.A (csr_minstret[63]), .Q
       (inc_ADD_UNS_OP_5_n_3782));
  INX1 inc_ADD_UNS_OP_5_g3490(.A (csr_minstret[60]), .Q
       (inc_ADD_UNS_OP_5_n_3785));
  INX1 inc_ADD_UNS_OP_5_g3492(.A (csr_minstret[41]), .Q
       (inc_ADD_UNS_OP_5_n_3789));
  INX1 inc_ADD_UNS_OP_5_g3493(.A (csr_minstret[44]), .Q
       (inc_ADD_UNS_OP_5_n_3791));
  INX1 inc_ADD_UNS_OP_5_g3494(.A (csr_minstret[62]), .Q
       (inc_ADD_UNS_OP_5_n_3792));
  INX1 inc_ADD_UNS_OP_5_g3495(.A (csr_minstret[54]), .Q
       (inc_ADD_UNS_OP_5_n_3793));
  INX1 inc_ADD_UNS_OP_5_g3496(.A (csr_minstret[56]), .Q
       (inc_ADD_UNS_OP_5_n_3795));
  INX1 inc_ADD_UNS_OP_5_g3497(.A (csr_minstret[38]), .Q
       (inc_ADD_UNS_OP_5_n_3798));
  INX1 inc_ADD_UNS_OP_5_g3498(.A (csr_minstret[43]), .Q
       (inc_ADD_UNS_OP_5_n_3800));
  INX1 inc_ADD_UNS_OP_5_g3500(.A (csr_minstret[58]), .Q
       (inc_ADD_UNS_OP_5_n_3803));
  INX1 inc_ADD_UNS_OP_5_g3502(.A (csr_minstret[42]), .Q
       (inc_ADD_UNS_OP_5_n_3808));
  INX1 inc_ADD_UNS_OP_5_g3504(.A (csr_minstret[39]), .Q
       (inc_ADD_UNS_OP_5_n_3812));
  INX1 inc_ADD_UNS_OP_5_g3506(.A (csr_minstret[40]), .Q
       (inc_ADD_UNS_OP_5_n_3815));
  INX1 inc_ADD_UNS_OP_5_g3510(.A (csr_minstret[51]), .Q
       (inc_ADD_UNS_OP_5_n_3824));
  INX1 inc_ADD_UNS_OP_5_g3511(.A (csr_minstret[49]), .Q
       (inc_ADD_UNS_OP_5_n_3826));
  INX1 inc_ADD_UNS_OP_5_g3514(.A (csr_minstret[53]), .Q
       (inc_ADD_UNS_OP_5_n_3832));
  INX1 inc_ADD_UNS_OP_5_g3515(.A (csr_minstret[32]), .Q
       (inc_ADD_UNS_OP_5_n_3834));
  INX1 inc_ADD_UNS_OP_5_g3517(.A (csr_minstret[47]), .Q
       (inc_ADD_UNS_OP_5_n_3838));
  EO2X1 inc_ADD_UNS_OP_5_g2(.A (inc_ADD_UNS_OP_5_n_3438), .B
       (csr_minstret[61]), .Q (n_7404));
  EO2X1 inc_ADD_UNS_OP_5_g3519(.A (inc_ADD_UNS_OP_5_n_3447), .B
       (csr_minstret[52]), .Q (n_7413));
  EO2X1 inc_ADD_UNS_OP_5_g3520(.A (inc_ADD_UNS_OP_5_n_3435), .B
       (n_7379), .Q (n_7438));
  EO2X1 inc_ADD_UNS_OP_5_g3521(.A (inc_ADD_UNS_OP_5_n_3476), .B
       (csr_minstret[59]), .Q (n_7406));
  EO2X1 inc_ADD_UNS_OP_5_g3522(.A (inc_ADD_UNS_OP_5_n_3474), .B
       (n_7381), .Q (n_7440));
  EO2X1 inc_ADD_UNS_OP_5_g3523(.A (inc_ADD_UNS_OP_5_n_3509), .B
       (csr_minstret[57]), .Q (n_7408));
  EO2X1 inc_ADD_UNS_OP_5_g3524(.A (inc_ADD_UNS_OP_5_n_3515), .B
       (csr_minstret[48]), .Q (n_7417));
  EO2X1 inc_ADD_UNS_OP_5_g3525(.A (inc_ADD_UNS_OP_5_n_3522), .B
       (n_7383), .Q (n_7442));
  EO2X1 inc_ADD_UNS_OP_5_g3526(.A (inc_ADD_UNS_OP_5_n_3536), .B
       (csr_minstret[46]), .Q (n_7419));
  EO2X1 inc_ADD_UNS_OP_5_g3527(.A (inc_ADD_UNS_OP_5_n_3580), .B
       (n_7387), .Q (n_7446));
  EO2X1 inc_ADD_UNS_OP_5_g3528(.A (inc_ADD_UNS_OP_5_n_3605), .B
       (n_7389), .Q (n_7448));
  MU2IX1 inc_ADD_UNS_OP_5_g3529(.S (inc_ADD_UNS_OP_5_n_3611), .IN0
       (inc_ADD_UNS_OP_5_n_3789), .IN1 (csr_minstret[41]), .Q (n_7424));
  EO2X1 inc_ADD_UNS_OP_5_g3530(.A (inc_ADD_UNS_OP_5_n_3621), .B
       (n_7391), .Q (n_7450));
  EO2X1 inc_ADD_UNS_OP_5_g3531(.A (inc_ADD_UNS_OP_5_n_3643), .B
       (n_7393), .Q (n_7452));
  EN2X1 inc_ADD_UNS_OP_5_g3532(.A (inc_ADD_UNS_OP_5_n_3681), .B
       (n_6232), .Q (n_7460));
  EO2X1 inc_ADD_UNS_OP_5_g3533(.A (inc_ADD_UNS_OP_5_n_3541), .B
       (n_7385), .Q (n_7444));
  EO2X1 inc_ADD_UNS_OP_5_g3534(.A (inc_ADD_UNS_OP_5_n_3655), .B
       (n_7395), .Q (n_7454));
  EN2X1 inc_ADD_UNS_OP_5_g3536(.A (inc_ADD_UNS_OP_5_n_3469), .B
       (csr_minstret[34]), .Q (n_7431));
  EO2X1 inc_ADD_UNS_OP_5_g3537(.A (inc_ADD_UNS_OP_5_n_3482), .B
       (csr_minstret[50]), .Q (n_7415));
  OR5X1 inc_ADD_UNS_OP_5_g3539(.A (inc_ADD_UNS_OP_5_n_3637), .B
       (inc_ADD_UNS_OP_5_n_3812), .C (inc_ADD_UNS_OP_5_n_3798), .D
       (inc_ADD_UNS_OP_5_n_3815), .E (inc_ADD_UNS_OP_5_n_3789), .Q
       (inc_ADD_UNS_OP_5_n_3597));
  MU2IX1 inc_add_1343_59_4_g3289(.S (inc_add_1343_59_4_n_3391), .IN0
       (csr_mcycle[32]), .IN1 (inc_add_1343_59_4_n_3786), .Q (n_7975));
  NO2X4 inc_add_1343_59_4_g3290(.A (inc_add_1343_59_4_n_3391), .B
       (inc_add_1343_59_4_n_3786), .Q (inc_add_1343_59_4_n_3386));
  NA2X4 inc_add_1343_59_4_g3292(.A (inc_add_1343_59_4_n_3403), .B
       (n_7635), .Q (inc_add_1343_59_4_n_3391));
  MU2IX1 inc_add_1343_59_4_g3297(.S (inc_add_1343_59_4_n_3419), .IN0
       (n_7376), .IN1 (inc_ADD_UNS_OP_5_n_3752), .Q (n_7977));
  NO2X4 inc_add_1343_59_4_g3299(.A (inc_add_1343_59_4_n_3419), .B
       (inc_ADD_UNS_OP_5_n_3752), .Q (inc_add_1343_59_4_n_3403));
  MU2IX1 inc_add_1343_59_4_g3302(.S (inc_add_1343_59_4_n_3428), .IN0
       (csr_mcycle[54]), .IN1 (inc_add_1343_59_4_n_3779), .Q (n_7921));
  NO2X2 inc_add_1343_59_4_g3303(.A (inc_add_1343_59_4_n_3428), .B
       (inc_add_1343_59_4_n_3779), .Q (inc_add_1343_59_4_n_3413));
  MU2IX1 inc_add_1343_59_4_g3305(.S (inc_add_1343_59_4_n_3440), .IN0
       (csr_mcycle[62]), .IN1 (inc_add_1343_59_4_n_3766), .Q (n_7913));
  NA2X4 inc_add_1343_59_4_g3306(.A (inc_add_1343_59_4_n_3435), .B
       (n_7377), .Q (inc_add_1343_59_4_n_3419));
  NO2X4 inc_add_1343_59_4_g3308(.A (inc_add_1343_59_4_n_3440), .B
       (inc_add_1343_59_4_n_3766), .Q (inc_add_1343_59_4_n_3423));
  NA2X4 inc_add_1343_59_4_g3310(.A (inc_add_1343_59_4_n_3432), .B
       (csr_mcycle[53]), .Q (inc_add_1343_59_4_n_3428));
  MU2IX1 inc_add_1343_59_4_g3311(.S (inc_add_1343_59_4_n_3446), .IN0
       (n_7378), .IN1 (inc_add_1345_58_1_n_3455), .Q (n_7979));
  HAX2 inc_add_1343_59_4_g3313(.A (inc_add_1343_59_4_n_3451), .B
       (csr_mcycle[52]), .S (n_7924), .CO (inc_add_1343_59_4_n_3432));
  NO2X4 inc_add_1343_59_4_g3316(.A (inc_add_1343_59_4_n_3446), .B
       (inc_add_1345_58_1_n_3455), .Q (inc_add_1343_59_4_n_3435));
  NA2X4 inc_add_1343_59_4_g3317(.A (inc_add_1343_59_4_n_3443), .B
       (csr_mcycle[61]), .Q (inc_add_1343_59_4_n_3440));
  HAX2 inc_add_1343_59_4_g3319(.A (inc_add_1343_59_4_n_3462), .B
       (csr_mcycle[60]), .S (n_7915), .CO (inc_add_1343_59_4_n_3443));
  NA2X4 inc_add_1343_59_4_g3321(.A (inc_add_1343_59_4_n_3457), .B
       (n_7379), .Q (inc_add_1343_59_4_n_3446));
  MU2IX1 inc_add_1343_59_4_g3323(.S (inc_add_1343_59_4_n_3468), .IN0
       (csr_mcycle[51]), .IN1 (inc_add_1343_59_4_n_3788), .Q (n_7928));
  NO2X4 inc_add_1343_59_4_g3324(.A (inc_add_1343_59_4_n_3468), .B
       (inc_add_1343_59_4_n_3788), .Q (inc_add_1343_59_4_n_3451));
  MU2IX1 inc_add_1343_59_4_g3325(.S (inc_add_1343_59_4_n_3475), .IN0
       (n_7380), .IN1 (inc_ADD_UNS_OP_5_n_3775), .Q (n_7981));
  MU2IX1 inc_add_1343_59_4_g3326(.S (inc_add_1343_59_4_n_3481), .IN0
       (csr_mcycle[59]), .IN1 (inc_add_1343_59_4_n_3758), .Q (n_7916));
  NO2X4 inc_add_1343_59_4_g3328(.A (inc_add_1343_59_4_n_3475), .B
       (inc_ADD_UNS_OP_5_n_3775), .Q (inc_add_1343_59_4_n_3457));
  NO2X4 inc_add_1343_59_4_g3329(.A (inc_add_1343_59_4_n_3481), .B
       (inc_add_1343_59_4_n_3758), .Q (inc_add_1343_59_4_n_3462));
  NA2X4 inc_add_1343_59_4_g3332(.A (inc_add_1343_59_4_n_3486), .B
       (csr_mcycle[50]), .Q (inc_add_1343_59_4_n_3468));
  NA2X4 inc_add_1343_59_4_g3337(.A (inc_add_1343_59_4_n_3492), .B
       (n_7381), .Q (inc_add_1343_59_4_n_3475));
  BUX1 inc_add_1343_59_4_g3339(.A (inc_add_1343_59_4_n_3492), .Q
       (inc_add_1343_59_4_n_3479));
  NA2X4 inc_add_1343_59_4_g3340(.A (inc_add_1343_59_4_n_3496), .B
       (csr_mcycle[58]), .Q (inc_add_1343_59_4_n_3481));
  MU2IX1 inc_add_1343_59_4_g3341(.S (inc_add_1343_59_4_n_3501), .IN0
       (csr_mcycle[49]), .IN1 (inc_add_1343_59_4_n_3784), .Q (n_7957));
  NO2X4 inc_add_1343_59_4_g3343(.A (inc_add_1343_59_4_n_3501), .B
       (inc_add_1343_59_4_n_3784), .Q (inc_add_1343_59_4_n_3486));
  MU2IX1 inc_add_1343_59_4_g3344(.S (inc_add_1343_59_4_n_3508), .IN0
       (n_8571), .IN1 (inc_ADD_UNS_OP_5_n_3756), .Q (n_7983));
  MU2IX1 inc_add_1343_59_4_g3345(.S (inc_add_1343_59_4_n_3512), .IN0
       (csr_mcycle[57]), .IN1 (inc_add_1343_59_4_n_3775), .Q (n_7918));
  NO2X4 inc_add_1343_59_4_g3346(.A (inc_add_1343_59_4_n_3508), .B
       (inc_ADD_UNS_OP_5_n_3756), .Q (inc_add_1343_59_4_n_3492));
  NO2X4 inc_add_1343_59_4_g3347(.A (inc_add_1343_59_4_n_3512), .B
       (inc_add_1343_59_4_n_3775), .Q (inc_add_1343_59_4_n_3496));
  NA2X4 inc_add_1343_59_4_g3349(.A (inc_add_1343_59_4_n_3505), .B
       (csr_mcycle[48]), .Q (inc_add_1343_59_4_n_3501));
  HAX2 inc_add_1343_59_4_g3352(.A (inc_add_1343_59_4_n_3524), .B
       (csr_mcycle[47]), .S (n_7959), .CO (inc_add_1343_59_4_n_3505));
  NA2X4 inc_add_1343_59_4_g3354(.A (inc_add_1343_59_4_n_3519), .B
       (n_7383), .Q (inc_add_1343_59_4_n_3508));
  NA2X4 inc_add_1343_59_4_g3356(.A (inc_add_1343_59_4_n_3805), .B
       (csr_mcycle[56]), .Q (inc_add_1343_59_4_n_3512));
  MU2IX1 inc_add_1343_59_4_g3359(.S (inc_add_1343_59_4_n_3527), .IN0
       (n_7384), .IN1 (inc_ADD_UNS_OP_5_n_3746), .Q (n_7985));
  NO2X4 inc_add_1343_59_4_g3361(.A (inc_add_1343_59_4_n_3527), .B
       (inc_ADD_UNS_OP_5_n_3746), .Q (inc_add_1343_59_4_n_3519));
  AND6X2 inc_add_1343_59_4_g3363(.A (inc_add_1343_59_4_n_3572), .B
       (csr_mcycle[42]), .C (csr_mcycle[44]), .D (csr_mcycle[43]), .E
       (csr_mcycle[45]), .F (csr_mcycle[46]), .Q
       (inc_add_1343_59_4_n_3524));
  NA2X4 inc_add_1343_59_4_g3365(.A (inc_add_1343_59_4_n_3539), .B
       (n_7385), .Q (inc_add_1343_59_4_n_3527));
  EO2X1 inc_add_1343_59_4_g3366(.A (inc_add_1343_59_4_n_3536), .B
       (csr_mcycle[45]), .Q (n_7961));
  NA2X1 inc_add_1343_59_4_g3367(.A (inc_add_1343_59_4_n_3536), .B
       (csr_mcycle[45]), .Q (inc_add_1343_59_4_n_3533));
  MU2IX1 inc_add_1343_59_4_g3368(.S (inc_add_1343_59_4_n_3544), .IN0
       (n_7386), .IN1 (inc_add_1343_59_4_n_3727), .Q (n_7987));
  HAX2 inc_add_1343_59_4_g3369(.A (inc_add_1343_59_4_n_3551), .B
       (csr_mcycle[44]), .S (n_7962), .CO (inc_add_1343_59_4_n_3536));
  NO2X4 inc_add_1343_59_4_g3370(.A (inc_add_1343_59_4_n_3544), .B
       (inc_add_1343_59_4_n_3727), .Q (inc_add_1343_59_4_n_3539));
  NA2X4 inc_add_1343_59_4_g3372(.A (inc_add_1343_59_4_n_3558), .B
       (n_7387), .Q (inc_add_1343_59_4_n_3544));
  EN2X1 inc_add_1343_59_4_g3373(.A (inc_add_1343_59_4_n_3806), .B
       (csr_mcycle[35]), .Q (n_7972));
  EO2X1 inc_add_1343_59_4_g3374(.A (inc_add_1343_59_4_n_3555), .B
       (csr_mcycle[43]), .Q (n_7963));
  AND5X1 inc_add_1343_59_4_g3375(.A (inc_add_1343_59_4_n_3583), .B
       (csr_mcycle[40]), .C (csr_mcycle[41]), .D (csr_mcycle[42]), .E
       (csr_mcycle[43]), .Q (inc_add_1343_59_4_n_3551));
  MU2IX1 inc_add_1343_59_4_g3376(.S (inc_add_1343_59_4_n_3561), .IN0
       (n_7388), .IN1 (inc_add_1343_59_4_n_3718), .Q (n_7989));
  HAX1 inc_add_1343_59_4_g3377(.A (inc_add_1343_59_4_n_3572), .B
       (csr_mcycle[42]), .S (n_7965), .CO (inc_add_1343_59_4_n_3555));
  NO2X4 inc_add_1343_59_4_g3379(.A (inc_add_1343_59_4_n_3561), .B
       (inc_add_1343_59_4_n_3718), .Q (inc_add_1343_59_4_n_3558));
  NA2X4 inc_add_1343_59_4_g3383(.A (inc_add_1343_59_4_n_3578), .B
       (n_7389), .Q (inc_add_1343_59_4_n_3561));
  EO2X1 inc_add_1343_59_4_g3384(.A (inc_add_1343_59_4_n_3576), .B
       (csr_mcycle[41]), .Q (n_7966));
  AND6X2 inc_add_1343_59_4_g3385(.A (inc_add_1343_59_4_n_3621), .B
       (csr_mcycle[37]), .C (csr_mcycle[39]), .D (csr_mcycle[38]), .E
       (csr_mcycle[40]), .F (csr_mcycle[41]), .Q
       (inc_add_1343_59_4_n_3572));
  HAX1 inc_add_1343_59_4_g3387(.A (inc_add_1343_59_4_n_3583), .B
       (csr_mcycle[40]), .S (n_7967), .CO (inc_add_1343_59_4_n_3576));
  NO2X4 inc_add_1343_59_4_g3388(.A (inc_add_1343_59_4_n_3586), .B
       (inc_add_1343_59_4_n_3736), .Q (inc_add_1343_59_4_n_3578));
  HAX1 inc_add_1343_59_4_g3391(.A (inc_add_1343_59_4_n_3592), .B
       (csr_mcycle[39]), .S (n_7968), .CO (inc_add_1343_59_4_n_3583));
  NA2X4 inc_add_1343_59_4_g3392(.A (inc_add_1343_59_4_n_3594), .B
       (n_7391), .Q (inc_add_1343_59_4_n_3586));
  HAX1 inc_add_1343_59_4_g3394(.A (inc_add_1343_59_4_n_3602), .B
       (csr_mcycle[38]), .S (n_7969), .CO (inc_add_1343_59_4_n_3592));
  NO2I1X4 inc_add_1343_59_4_g3395(.B (inc_add_1343_59_4_n_3605), .AN
       (n_7392), .Q (inc_add_1343_59_4_n_3594));
  EO2X1 inc_add_1343_59_4_g3398(.A (inc_add_1343_59_4_n_3614), .B
       (n_7393), .Q (n_7994));
  HAX1 inc_add_1343_59_4_g3399(.A (inc_add_1343_59_4_n_3621), .B
       (csr_mcycle[37]), .S (n_7970), .CO (inc_add_1343_59_4_n_3602));
  NA2X4 inc_add_1343_59_4_g3400(.A (inc_add_1343_59_4_n_3614), .B
       (n_7393), .Q (inc_add_1343_59_4_n_3605));
  EO2X1 inc_add_1343_59_4_g3401(.A (inc_add_1343_59_4_n_3611), .B
       (n_7399), .Q (n_8000));
  HAX1 inc_add_1343_59_4_g3402(.A (inc_add_1343_59_4_n_3620), .B
       (n_7400), .S (n_8001), .CO (inc_add_1343_59_4_n_3611));
  NO2I1X4 inc_add_1343_59_4_g3404(.B (inc_add_1343_59_4_n_3624), .AN
       (n_7394), .Q (inc_add_1343_59_4_n_3614));
  HAX1 inc_add_1343_59_4_g3407(.A (inc_add_1343_59_4_n_3633), .B
       (n_7401), .S (n_8002), .CO (inc_add_1343_59_4_n_3620));
  NO2I1X4 inc_add_1343_59_4_g3408(.B (inc_add_1343_59_4_n_3628), .AN
       (csr_mcycle[36]), .Q (inc_add_1343_59_4_n_3621));
  EO2X1 inc_add_1343_59_4_g3409(.A (inc_add_1343_59_4_n_3629), .B
       (n_7395), .Q (n_7996));
  NA2X4 inc_add_1343_59_4_g3410(.A (inc_add_1343_59_4_n_3635), .B
       (n_7395), .Q (inc_add_1343_59_4_n_3624));
  NA2X4 inc_add_1343_59_4_g3412(.A (inc_add_1343_59_4_n_3629), .B
       (inc_add_1343_59_4_n_3646), .Q (inc_add_1343_59_4_n_3628));
  BUX1 inc_add_1343_59_4_g3414(.A (inc_add_1343_59_4_n_3635), .Q
       (inc_add_1343_59_4_n_3629));
  HAX1 inc_add_1343_59_4_g3415(.A (inc_add_1343_59_4_n_3640), .B
       (n_7632), .S (n_8003), .CO (inc_add_1343_59_4_n_3633));
  NO2I1X4 inc_add_1343_59_4_g3417(.B (inc_add_1343_59_4_n_3642), .AN
       (n_8354), .Q (inc_add_1343_59_4_n_3635));
  HAX1 inc_add_1343_59_4_g3419(.A (inc_add_1343_59_4_n_3648), .B
       (n_8208), .S (n_8004), .CO (inc_add_1343_59_4_n_3640));
  EO2X1 inc_add_1343_59_4_g3420(.A (inc_add_1343_59_4_n_3653), .B
       (n_7397), .Q (n_7998));
  NA2X4 inc_add_1343_59_4_g3421(.A (inc_add_1343_59_4_n_3653), .B
       (n_7397), .Q (inc_add_1343_59_4_n_3642));
  NO3X4 inc_add_1343_59_4_g3422(.A (inc_add_1343_59_4_n_3656), .B
       (inc_add_1343_59_4_n_3658), .C (inc_add_1343_59_4_n_3663), .Q
       (inc_add_1343_59_4_n_3646));
  HAX1 inc_add_1343_59_4_g3423(.A (inc_add_1343_59_4_n_3696), .B
       (n_7633), .S (n_8005), .CO (inc_add_1343_59_4_n_3648));
  NO2X1 inc_add_1343_59_4_g3424(.A (inc_add_1343_59_4_n_3656), .B
       (inc_add_1343_59_4_n_3658), .Q (inc_add_1343_59_4_n_3649));
  EN2X0 inc_add_1343_59_4_g3425(.A (inc_add_1343_59_4_n_3664), .B
       (n_7398), .Q (n_7999));
  NO2I1X4 inc_add_1343_59_4_g3426(.B (inc_add_1343_59_4_n_3664), .AN
       (n_7398), .Q (inc_add_1343_59_4_n_3653));
  NA2X2 inc_add_1343_59_4_g3428(.A (inc_add_1343_59_4_n_3660), .B
       (inc_add_1343_59_4_n_3684), .Q (inc_add_1343_59_4_n_3656));
  NA3X2 inc_add_1343_59_4_g3429(.A (inc_add_1343_59_4_n_3687), .B
       (inc_add_1343_59_4_n_3681), .C (n_7384), .Q
       (inc_add_1343_59_4_n_3658));
  AND6X2 inc_add_1343_59_4_g3430(.A (n_7380), .B (n_7379), .C (n_7635),
       .D (n_7381), .E (csr_mcycle[32]), .F (csr_mcycle[33]), .Q
       (inc_add_1343_59_4_n_3660));
  NA2X2 inc_add_1343_59_4_g3431(.A (inc_add_1343_59_4_n_3680), .B
       (inc_add_1343_59_4_n_3674), .Q (inc_add_1343_59_4_n_3663));
  NA2X4 inc_add_1343_59_4_g3432(.A (inc_add_1343_59_4_n_3669), .B
       (inc_add_1343_59_4_n_3693), .Q (inc_add_1343_59_4_n_3664));
  NA5X1 inc_add_1343_59_4_g3433(.A (inc_add_1343_59_4_n_3677), .B
       (csr_mcycle[47]), .C (csr_mcycle[48]), .D (csr_mcycle[54]), .E
       (csr_mcycle[51]), .Q (inc_add_1343_59_4_n_3665));
  AND6X2 inc_add_1343_59_4_g3434(.A (n_7633), .B (n_7632), .C (n_8208),
       .D (n_7636), .E (n_6235), .F (n_7401), .Q
       (inc_add_1343_59_4_n_3669));
  AND5X2 inc_add_1343_59_4_g3435(.A (n_7395), .B (n_7394), .C (n_8622),
       .D (n_7389), .E (csr_mcycle[35]), .Q (inc_add_1343_59_4_n_3674));
  AND5X1 inc_add_1343_59_4_g3436(.A (csr_mcycle[49]), .B
       (csr_mcycle[55]), .C (csr_mcycle[50]), .D (csr_mcycle[52]), .E
       (csr_mcycle[53]), .Q (inc_add_1343_59_4_n_3677));
  AND3X1 inc_add_1343_59_4_g3437(.A (n_7392), .B (n_7391), .C (n_7393),
       .Q (inc_add_1343_59_4_n_3680));
  AND4X2 inc_add_1343_59_4_g3438(.A (n_7385), .B (n_7387), .C (n_8571),
       .D (n_7386), .Q (inc_add_1343_59_4_n_3681));
  AND3X1 inc_add_1343_59_4_g3439(.A (n_7376), .B (n_7378), .C (n_7377),
       .Q (inc_add_1343_59_4_n_3684));
  AND3X1 inc_add_1343_59_4_g3440(.A (n_7383), .B (n_7388), .C
       (csr_mcycle[34]), .Q (inc_add_1343_59_4_n_3687));
  EO2X1 inc_add_1343_59_4_g3441(.A (n_6235), .B (n_7636), .Q (n_8006));
  AND2X4 inc_add_1343_59_4_g3442(.A (n_7400), .B (n_7399), .Q
       (inc_add_1343_59_4_n_3693));
  AND2X1 inc_add_1343_59_4_g3443(.A (n_7636), .B (n_6235), .Q
       (inc_add_1343_59_4_n_3696));
  INX1 inc_add_1343_59_4_g3447(.A (n_7378), .Q
       (inc_add_1345_58_1_n_3455));
  INX1 inc_add_1343_59_4_g3450(.A (n_7388), .Q
       (inc_add_1343_59_4_n_3718));
  INX1 inc_add_1343_59_4_g3454(.A (n_7386), .Q
       (inc_add_1343_59_4_n_3727));
  INX1 inc_add_1343_59_4_g3458(.A (n_8622), .Q
       (inc_add_1343_59_4_n_3736));
  INX1 inc_add_1343_59_4_g3463(.A (csr_mcycle[55]), .Q
       (inc_add_1343_59_4_n_3749));
  INX1 inc_add_1343_59_4_g3466(.A (csr_mcycle[59]), .Q
       (inc_add_1343_59_4_n_3758));
  INX1 inc_add_1343_59_4_g3469(.A (csr_mcycle[62]), .Q
       (inc_add_1343_59_4_n_3766));
  INX1 inc_add_1343_59_4_g3470(.A (csr_mcycle[33]), .Q
       (inc_add_1343_59_4_n_3769));
  INX1 inc_add_1343_59_4_g3471(.A (csr_mcycle[57]), .Q
       (inc_add_1343_59_4_n_3775));
  INX1 inc_add_1343_59_4_g3472(.A (csr_mcycle[54]), .Q
       (inc_add_1343_59_4_n_3779));
  INX1 inc_add_1343_59_4_g3474(.A (csr_mcycle[49]), .Q
       (inc_add_1343_59_4_n_3784));
  INX1 inc_add_1343_59_4_g3475(.A (csr_mcycle[32]), .Q
       (inc_add_1343_59_4_n_3786));
  INX1 inc_add_1343_59_4_g3476(.A (csr_mcycle[51]), .Q
       (inc_add_1343_59_4_n_3788));
  EO2X1 inc_add_1343_59_4_g2(.A (inc_add_1343_59_4_n_3403), .B
       (n_7635), .Q (n_7976));
  EO2X1 inc_add_1343_59_4_g3479(.A (inc_add_1343_59_4_n_3435), .B
       (n_7377), .Q (n_7978));
  EO2X1 inc_add_1343_59_4_g3480(.A (inc_add_1343_59_4_n_3432), .B
       (csr_mcycle[53]), .Q (n_7922));
  EO2X1 inc_add_1343_59_4_g3481(.A (inc_add_1343_59_4_n_3443), .B
       (csr_mcycle[61]), .Q (n_7914));
  EO2X1 inc_add_1343_59_4_g3482(.A (inc_add_1343_59_4_n_3457), .B
       (n_7379), .Q (n_7980));
  EO2X1 inc_add_1343_59_4_g3483(.A (inc_add_1343_59_4_n_3486), .B
       (csr_mcycle[50]), .Q (n_7949));
  EO2X1 inc_add_1343_59_4_g3484(.A (inc_add_1343_59_4_n_3479), .B
       (n_7381), .Q (n_7982));
  EO2X1 inc_add_1343_59_4_g3485(.A (inc_add_1343_59_4_n_3496), .B
       (csr_mcycle[58]), .Q (n_7917));
  EO2X1 inc_add_1343_59_4_g3486(.A (inc_add_1343_59_4_n_3505), .B
       (csr_mcycle[48]), .Q (n_7958));
  EO2X1 inc_add_1343_59_4_g3487(.A (inc_add_1343_59_4_n_3519), .B
       (n_7383), .Q (n_7984));
  EO2X1 inc_add_1343_59_4_g3488(.A (inc_add_1343_59_4_n_3805), .B
       (csr_mcycle[56]), .Q (n_7919));
  NO2I1X4 inc_add_1343_59_4_g3489(.B (inc_add_1343_59_4_n_3665), .AN
       (inc_add_1343_59_4_n_3524), .Q (inc_add_1343_59_4_n_3805));
  NA2I1X1 inc_add_1343_59_4_g3490(.B (inc_add_1343_59_4_n_3649), .AN
       (inc_add_1343_59_4_n_3561), .Q (inc_add_1343_59_4_n_3806));
  MU2IX1 inc_add_1343_59_4_g3491(.S (inc_add_1343_59_4_n_3586), .IN0
       (n_8622), .IN1 (inc_add_1343_59_4_n_3736), .Q (n_7991));
  EN2X1 inc_add_1343_59_4_g3492(.A (n_7392), .B
       (inc_add_1343_59_4_n_3605), .Q (n_7993));
  EN2X1 inc_add_1343_59_4_g3493(.A (inc_add_1343_59_4_n_3624), .B
       (n_7394), .Q (n_7995));
  EN2X1 inc_add_1343_59_4_g3494(.A (inc_add_1343_59_4_n_3628), .B
       (csr_mcycle[36]), .Q (n_7971));
  EN2X1 inc_add_1343_59_4_g3495(.A (inc_add_1343_59_4_n_3642), .B
       (n_8354), .Q (n_7997));
  NA2I1X1 inc_add_1343_59_4_g3496(.B (inc_add_1343_59_4_n_3479), .AN
       (inc_add_1343_59_4_n_3656), .Q (inc_add_1343_59_4_n_3812));
  EO2X1 inc_add_1343_59_4_g3497(.A (inc_add_1343_59_4_n_3594), .B
       (n_7391), .Q (n_7992));
  EO2X1 inc_add_1343_59_4_g3498(.A (inc_add_1343_59_4_n_3558), .B
       (n_7387), .Q (n_7988));
  EO2X1 inc_add_1343_59_4_g3499(.A (inc_add_1343_59_4_n_3539), .B
       (n_7385), .Q (n_7986));
  EO2X1 inc_add_1343_59_4_g3500(.A (inc_add_1343_59_4_n_3578), .B
       (n_7389), .Q (n_7990));
  EN2X1 inc_add_1343_59_4_g3501(.A (inc_add_1343_59_4_n_3533), .B
       (csr_mcycle[46]), .Q (n_7960));
  EN2X1 inc_add_1343_59_4_g3502(.A (inc_add_1343_59_4_n_3812), .B
       (csr_mcycle[34]), .Q (n_7973));
  NA2X2 inc_ADD_UNS_OP5491_6_g2395(.A (inc_ADD_UNS_OP5491_6_n_2356), .B
       (n_7376), .Q (inc_ADD_UNS_OP5491_6_n_2351));
  MU2IX1 inc_ADD_UNS_OP5491_6_g2397(.S (inc_ADD_UNS_OP5491_6_n_2362),
       .IN0 (n_7377), .IN1 (inc_ADD_UNS_OP5491_6_n_2657), .Q (n_7471));
  NO2X4 inc_ADD_UNS_OP5491_6_g2398(.A (inc_ADD_UNS_OP5491_6_n_2362), .B
       (inc_ADD_UNS_OP5491_6_n_2657), .Q (inc_ADD_UNS_OP5491_6_n_2356));
  NA2X2 inc_ADD_UNS_OP5491_6_g2401(.A (inc_ADD_UNS_OP5491_6_n_2366), .B
       (n_7378), .Q (inc_ADD_UNS_OP5491_6_n_2362));
  MU2IX1 inc_ADD_UNS_OP5491_6_g2404(.S (inc_ADD_UNS_OP5491_6_n_2372),
       .IN0 (n_7379), .IN1 (inc_ADD_UNS_OP5491_6_n_2641), .Q (n_7475));
  NO2X4 inc_ADD_UNS_OP5491_6_g2405(.A (inc_ADD_UNS_OP5491_6_n_2372), .B
       (inc_ADD_UNS_OP5491_6_n_2641), .Q (inc_ADD_UNS_OP5491_6_n_2366));
  NA2X2 inc_ADD_UNS_OP5491_6_g2408(.A (inc_ADD_UNS_OP5491_6_n_2380), .B
       (n_7380), .Q (inc_ADD_UNS_OP5491_6_n_2372));
  AND6X2 inc_ADD_UNS_OP5491_6_g2411(.A (inc_ADD_UNS_OP5491_6_n_2410),
       .B (n_7384), .C (n_7385), .D (n_7383), .E (n_8571), .F (n_7381),
       .Q (inc_ADD_UNS_OP5491_6_n_2380));
  NA2X1 inc_ADD_UNS_OP5491_6_g2415(.A (inc_ADD_UNS_OP5491_6_n_2393), .B
       (n_8571), .Q (inc_ADD_UNS_OP5491_6_n_2388));
  MU2IX1 inc_ADD_UNS_OP5491_6_g2417(.S (inc_ADD_UNS_OP5491_6_n_2399),
       .IN0 (n_7383), .IN1 (n_8655), .Q (n_7483));
  NO2X1 inc_ADD_UNS_OP5491_6_g2418(.A (inc_ADD_UNS_OP5491_6_n_2399), .B
       (n_8655), .Q (inc_ADD_UNS_OP5491_6_n_2393));
  NA2X1 inc_ADD_UNS_OP5491_6_g2420(.A (inc_ADD_UNS_OP5491_6_n_2401), .B
       (n_7384), .Q (inc_ADD_UNS_OP5491_6_n_2399));
  AND6X2 inc_ADD_UNS_OP5491_6_g2423(.A (inc_ADD_UNS_OP5491_6_n_2431),
       .B (n_7387), .C (n_7388), .D (n_7386), .E (n_7385), .F (n_7389),
       .Q (inc_ADD_UNS_OP5491_6_n_2401));
  AND6X2 inc_ADD_UNS_OP5491_6_g2426(.A (inc_ADD_UNS_OP5491_6_n_2438),
       .B (n_7388), .C (n_7387), .D (n_7386), .E (n_8622), .F (n_7389),
       .Q (inc_ADD_UNS_OP5491_6_n_2410));
  NA2X1 inc_ADD_UNS_OP5491_6_g2430(.A (inc_ADD_UNS_OP5491_6_n_2421), .B
       (n_7387), .Q (inc_ADD_UNS_OP5491_6_n_2419));
  HAX2 inc_ADD_UNS_OP5491_6_g2432(.A (inc_ADD_UNS_OP5491_6_n_2424), .B
       (n_7388), .S (n_7493), .CO (inc_ADD_UNS_OP5491_6_n_2421));
  AND6X2 inc_ADD_UNS_OP5491_6_g2434(.A (inc_ADD_UNS_OP5491_6_n_2460),
       .B (n_7392), .C (n_7391), .D (n_7393), .E (n_8622), .F (n_7389),
       .Q (inc_ADD_UNS_OP5491_6_n_2424));
  AND6X2 inc_ADD_UNS_OP5491_6_g2438(.A (inc_ADD_UNS_OP5491_6_n_2468),
       .B (n_7392), .C (n_7394), .D (n_7391), .E (n_7393), .F (n_8622),
       .Q (inc_ADD_UNS_OP5491_6_n_2431));
  AND6X2 inc_ADD_UNS_OP5491_6_g2441(.A (inc_ADD_UNS_OP5491_6_n_2476),
       .B (n_7392), .C (n_7395), .D (n_7393), .E (n_7394), .F (n_7391),
       .Q (inc_ADD_UNS_OP5491_6_n_2438));
  NA2X1 inc_ADD_UNS_OP5491_6_g2442(.A (inc_ADD_UNS_OP5491_6_n_2443), .B
       (n_6233), .Q (inc_ADD_UNS_OP5491_6_n_2440));
  HAX2 inc_ADD_UNS_OP5491_6_g2443(.A (inc_ADD_UNS_OP5491_6_n_2450), .B
       (n_6235), .S (n_7527), .CO (inc_ADD_UNS_OP5491_6_n_2443));
  NA2X1 inc_ADD_UNS_OP5491_6_g2445(.A (inc_ADD_UNS_OP5491_6_n_2452), .B
       (n_7392), .Q (inc_ADD_UNS_OP5491_6_n_2446));
  HAX2 inc_ADD_UNS_OP5491_6_g2447(.A (inc_ADD_UNS_OP5491_6_n_2458), .B
       (n_6236), .S (n_7529), .CO (inc_ADD_UNS_OP5491_6_n_2450));
  MU2IX1 inc_ADD_UNS_OP5491_6_g2448(.S (inc_ADD_UNS_OP5491_6_n_2455),
       .IN0 (n_7393), .IN1 (inc_ADD_UNS_OP5491_6_n_2675), .Q (n_7503));
  NO2X1 inc_ADD_UNS_OP5491_6_g2449(.A (inc_ADD_UNS_OP5491_6_n_2455), .B
       (inc_ADD_UNS_OP5491_6_n_2675), .Q (inc_ADD_UNS_OP5491_6_n_2452));
  INX1 inc_ADD_UNS_OP5491_6_g2450(.A (inc_ADD_UNS_OP5491_6_n_2460), .Q
       (inc_ADD_UNS_OP5491_6_n_2455));
  HAX2 inc_ADD_UNS_OP5491_6_g2451(.A (inc_ADD_UNS_OP5491_6_n_2463), .B
       (csr_minstret[31]), .S (n_7531), .CO
       (inc_ADD_UNS_OP5491_6_n_2458));
  HAX2 inc_ADD_UNS_OP5491_6_g2454(.A (inc_ADD_UNS_OP5491_6_n_2473), .B
       (csr_minstret[30]), .S (n_7533), .CO
       (inc_ADD_UNS_OP5491_6_n_2463));
  AND6X2 inc_ADD_UNS_OP5491_6_g2457(.A (inc_ADD_UNS_OP5491_6_n_2503),
       .B (n_6238), .C (n_8354), .D (n_7395), .E (n_7398), .F (n_7397),
       .Q (inc_ADD_UNS_OP5491_6_n_2468));
  HAX2 inc_ADD_UNS_OP5491_6_g2458(.A (inc_ADD_UNS_OP5491_6_n_2481), .B
       (csr_minstret[29]), .S (n_7535), .CO
       (inc_ADD_UNS_OP5491_6_n_2473));
  EO2X1 inc_ADD_UNS_OP5491_6_g2459(.A (inc_ADD_UNS_OP5491_6_n_2479), .B
       (n_8354), .Q (n_7509));
  AND6X2 inc_ADD_UNS_OP5491_6_g2460(.A (inc_ADD_UNS_OP5491_6_n_2515),
       .B (n_6237), .C (n_6238), .D (n_8354), .E (n_7398), .F (n_7397),
       .Q (inc_ADD_UNS_OP5491_6_n_2476));
  HAX1 inc_ADD_UNS_OP5491_6_g2461(.A (inc_ADD_UNS_OP5491_6_n_2484), .B
       (n_7397), .S (n_7511), .CO (inc_ADD_UNS_OP5491_6_n_2479));
  HAX1 inc_ADD_UNS_OP5491_6_g2464(.A (inc_ADD_UNS_OP5491_6_n_2497), .B
       (n_7398), .S (n_7513), .CO (inc_ADD_UNS_OP5491_6_n_2484));
  EO2X1 inc_ADD_UNS_OP5491_6_g2466(.A (inc_ADD_UNS_OP5491_6_n_2493), .B
       (csr_minstret[27]), .Q (n_7539));
  NA2X1 inc_ADD_UNS_OP5491_6_g2467(.A (inc_ADD_UNS_OP5491_6_n_2493), .B
       (csr_minstret[27]), .Q (inc_ADD_UNS_OP5491_6_n_2489));
  HAX2 inc_ADD_UNS_OP5491_6_g2468(.A (inc_ADD_UNS_OP5491_6_n_2507), .B
       (csr_minstret[26]), .S (n_7541), .CO
       (inc_ADD_UNS_OP5491_6_n_2493));
  EO2X1 inc_ADD_UNS_OP5491_6_g2469(.A (inc_ADD_UNS_OP5491_6_n_2503), .B
       (n_6238), .Q (n_7515));
  AND5X1 inc_ADD_UNS_OP5491_6_g2470(.A (inc_ADD_UNS_OP5491_6_n_2526),
       .B (inc_ADD_UNS_OP5491_6_n_2611), .C (n_6237), .D (n_6238), .E
       (n_6232), .Q (inc_ADD_UNS_OP5491_6_n_2497));
  EO2X1 inc_ADD_UNS_OP5491_6_g2471(.A (inc_ADD_UNS_OP5491_6_n_2515), .B
       (n_6237), .Q (n_7517));
  AND6X2 inc_ADD_UNS_OP5491_6_g2473(.A (inc_ADD_UNS_OP5491_6_n_2531),
       .B (inc_ADD_UNS_OP5491_6_n_2611), .C (n_6233), .D (n_6237), .E
       (n_6234), .F (n_6232), .Q (inc_ADD_UNS_OP5491_6_n_2503));
  EO2X1 inc_ADD_UNS_OP5491_6_g2476(.A (inc_ADD_UNS_OP5491_6_n_2521), .B
       (n_7632), .Q (n_7521));
  EN2X0 inc_ADD_UNS_OP5491_6_g2477(.A (inc_ADD_UNS_OP5491_6_n_2523), .B
       (n_6232), .Q (n_7519));
  EO2X1 inc_ADD_UNS_OP5491_6_g2478(.A (inc_ADD_UNS_OP5491_6_n_2527), .B
       (csr_minstret[24]), .Q (n_7545));
  NO2I1X2 inc_ADD_UNS_OP5491_6_g2479(.B (inc_ADD_UNS_OP5491_6_n_2523),
       .AN (n_6232), .Q (inc_ADD_UNS_OP5491_6_n_2515));
  NA2X2 inc_ADD_UNS_OP5491_6_g2480(.A (inc_ADD_UNS_OP5491_6_n_2527), .B
       (csr_minstret[24]), .Q (inc_ADD_UNS_OP5491_6_n_2517));
  NO2I1X1 inc_ADD_UNS_OP5491_6_g2481(.B (inc_ADD_UNS_OP5491_6_n_2616),
       .AN (inc_ADD_UNS_OP5491_6_n_2526), .Q
       (inc_ADD_UNS_OP5491_6_n_2521));
  NA2X1 inc_ADD_UNS_OP5491_6_g2482(.A (inc_ADD_UNS_OP5491_6_n_2526), .B
       (inc_ADD_UNS_OP5491_6_n_2611), .Q (inc_ADD_UNS_OP5491_6_n_2523));
  EO2X1 inc_ADD_UNS_OP5491_6_g2483(.A (inc_ADD_UNS_OP5491_6_n_2531), .B
       (csr_minstret[23]), .Q (n_7547));
  AND3X2 inc_ADD_UNS_OP5491_6_g2484(.A (inc_ADD_UNS_OP5491_6_n_2531),
       .B (n_6233), .C (n_6234), .Q (inc_ADD_UNS_OP5491_6_n_2526));
  AND2X4 inc_ADD_UNS_OP5491_6_g2485(.A (inc_ADD_UNS_OP5491_6_n_2531),
       .B (csr_minstret[23]), .Q (inc_ADD_UNS_OP5491_6_n_2527));
  EO2X1 inc_ADD_UNS_OP5491_6_g2486(.A (inc_ADD_UNS_OP5491_6_n_2534), .B
       (csr_minstret[22]), .Q (n_7549));
  AND5X2 inc_ADD_UNS_OP5491_6_g2487(.A (inc_ADD_UNS_OP5491_6_n_2543),
       .B (csr_minstret[19]), .C (csr_minstret[20]), .D
       (csr_minstret[21]), .E (csr_minstret[22]), .Q
       (inc_ADD_UNS_OP5491_6_n_2531));
  HAX1 inc_ADD_UNS_OP5491_6_g2488(.A (inc_ADD_UNS_OP5491_6_n_2537), .B
       (csr_minstret[21]), .S (n_7551), .CO
       (inc_ADD_UNS_OP5491_6_n_2534));
  HAX1 inc_ADD_UNS_OP5491_6_g2489(.A (inc_ADD_UNS_OP5491_6_n_2540), .B
       (csr_minstret[20]), .S (n_7553), .CO
       (inc_ADD_UNS_OP5491_6_n_2537));
  HAX1 inc_ADD_UNS_OP5491_6_g2490(.A (inc_ADD_UNS_OP5491_6_n_2543), .B
       (csr_minstret[19]), .S (n_7555), .CO
       (inc_ADD_UNS_OP5491_6_n_2540));
  HAX1 inc_ADD_UNS_OP5491_6_g2491(.A (inc_ADD_UNS_OP5491_6_n_2546), .B
       (csr_minstret[18]), .S (n_7557), .CO
       (inc_ADD_UNS_OP5491_6_n_2543));
  HAX1 inc_ADD_UNS_OP5491_6_g2492(.A (inc_ADD_UNS_OP5491_6_n_2548), .B
       (csr_minstret[17]), .S (n_7559), .CO
       (inc_ADD_UNS_OP5491_6_n_2546));
  EO2X1 inc_ADD_UNS_OP5491_6_g2493(.A (inc_ADD_UNS_OP5491_6_n_2551), .B
       (csr_minstret[16]), .Q (n_7561));
  AND3X2 inc_ADD_UNS_OP5491_6_g2494(.A (inc_ADD_UNS_OP5491_6_n_2556),
       .B (csr_minstret[15]), .C (csr_minstret[16]), .Q
       (inc_ADD_UNS_OP5491_6_n_2548));
  HAX1 inc_ADD_UNS_OP5491_6_g2495(.A (inc_ADD_UNS_OP5491_6_n_2556), .B
       (csr_minstret[15]), .S (n_7563), .CO
       (inc_ADD_UNS_OP5491_6_n_2551));
  EO2X0 inc_ADD_UNS_OP5491_6_g2496(.A (inc_ADD_UNS_OP5491_6_n_2561), .B
       (csr_minstret[14]), .Q (n_7565));
  AND2X2 inc_ADD_UNS_OP5491_6_g2497(.A (inc_ADD_UNS_OP5491_6_n_2561),
       .B (csr_minstret[14]), .Q (inc_ADD_UNS_OP5491_6_n_2556));
  EO2X0 inc_ADD_UNS_OP5491_6_g2498(.A (inc_ADD_UNS_OP5491_6_n_2566), .B
       (csr_minstret[13]), .Q (n_7567));
  AND2X2 inc_ADD_UNS_OP5491_6_g2499(.A (inc_ADD_UNS_OP5491_6_n_2566),
       .B (csr_minstret[13]), .Q (inc_ADD_UNS_OP5491_6_n_2561));
  EO2X0 inc_ADD_UNS_OP5491_6_g2500(.A (inc_ADD_UNS_OP5491_6_n_2571), .B
       (csr_minstret[12]), .Q (n_7569));
  AND2X1 inc_ADD_UNS_OP5491_6_g2501(.A (inc_ADD_UNS_OP5491_6_n_2571),
       .B (csr_minstret[12]), .Q (inc_ADD_UNS_OP5491_6_n_2566));
  EO2X0 inc_ADD_UNS_OP5491_6_g2502(.A (inc_ADD_UNS_OP5491_6_n_2576), .B
       (csr_minstret[11]), .Q (n_7571));
  AND2X1 inc_ADD_UNS_OP5491_6_g2503(.A (inc_ADD_UNS_OP5491_6_n_2576),
       .B (csr_minstret[11]), .Q (inc_ADD_UNS_OP5491_6_n_2571));
  EO2X1 inc_ADD_UNS_OP5491_6_g2504(.A (inc_ADD_UNS_OP5491_6_n_2581), .B
       (csr_minstret[10]), .Q (n_7573));
  AND2X2 inc_ADD_UNS_OP5491_6_g2505(.A (inc_ADD_UNS_OP5491_6_n_2581),
       .B (csr_minstret[10]), .Q (inc_ADD_UNS_OP5491_6_n_2576));
  EO2X0 inc_ADD_UNS_OP5491_6_g2506(.A (inc_ADD_UNS_OP5491_6_n_2586), .B
       (csr_minstret[9]), .Q (n_7575));
  AND2X4 inc_ADD_UNS_OP5491_6_g2507(.A (inc_ADD_UNS_OP5491_6_n_2586),
       .B (csr_minstret[9]), .Q (inc_ADD_UNS_OP5491_6_n_2581));
  EO2X0 inc_ADD_UNS_OP5491_6_g2508(.A (inc_ADD_UNS_OP5491_6_n_2591), .B
       (csr_minstret[8]), .Q (n_7577));
  AND2X4 inc_ADD_UNS_OP5491_6_g2509(.A (inc_ADD_UNS_OP5491_6_n_2591),
       .B (csr_minstret[8]), .Q (inc_ADD_UNS_OP5491_6_n_2586));
  NO2I1X2 inc_ADD_UNS_OP5491_6_g2511(.B (inc_ADD_UNS_OP5491_6_n_2596),
       .AN (csr_minstret[7]), .Q (inc_ADD_UNS_OP5491_6_n_2591));
  EO2X0 inc_ADD_UNS_OP5491_6_g2513(.A (inc_ADD_UNS_OP5491_6_n_2601), .B
       (csr_minstret[6]), .Q (n_7581));
  NA2X2 inc_ADD_UNS_OP5491_6_g2514(.A (inc_ADD_UNS_OP5491_6_n_2601), .B
       (csr_minstret[6]), .Q (inc_ADD_UNS_OP5491_6_n_2596));
  EO2X0 inc_ADD_UNS_OP5491_6_g2515(.A (inc_ADD_UNS_OP5491_6_n_2606), .B
       (csr_minstret[5]), .Q (n_7583));
  AND2X4 inc_ADD_UNS_OP5491_6_g2516(.A (inc_ADD_UNS_OP5491_6_n_2606),
       .B (csr_minstret[5]), .Q (inc_ADD_UNS_OP5491_6_n_2601));
  NO2I1X2 inc_ADD_UNS_OP5491_6_g2518(.B (inc_ADD_UNS_OP5491_6_n_2620),
       .AN (csr_minstret[4]), .Q (inc_ADD_UNS_OP5491_6_n_2606));
  EO2X1 inc_ADD_UNS_OP5491_6_g2519(.A (inc_ADD_UNS_OP5491_6_n_2615), .B
       (csr_minstret[2]), .Q (n_7589));
  NO2I1X1 inc_ADD_UNS_OP5491_6_g2521(.B (inc_ADD_UNS_OP5491_6_n_2616),
       .AN (n_7632), .Q (inc_ADD_UNS_OP5491_6_n_2611));
  HAX1 inc_ADD_UNS_OP5491_6_g2522(.A (inc_ADD_UNS_OP5491_6_n_2626), .B
       (csr_minstret[1]), .S (n_7591), .CO
       (inc_ADD_UNS_OP5491_6_n_2615));
  NA3X1 inc_ADD_UNS_OP5491_6_g2523(.A (n_6236), .B (n_6235), .C
       (inc_ADD_UNS_OP5491_6_n_2622), .Q (inc_ADD_UNS_OP5491_6_n_2616));
  NA2X2 inc_ADD_UNS_OP5491_6_g2525(.A (inc_ADD_UNS_OP5491_6_n_2625), .B
       (csr_minstret[3]), .Q (inc_ADD_UNS_OP5491_6_n_2620));
  AND6X1 inc_ADD_UNS_OP5491_6_g2526(.A (inc_ADD_UNS_OP5491_6_n_2628),
       .B (csr_minstret[27]), .C (csr_minstret[25]), .D
       (csr_minstret[24]), .E (csr_minstret[26]), .F
       (csr_minstret[23]), .Q (inc_ADD_UNS_OP5491_6_n_2622));
  NO2X2 inc_ADD_UNS_OP5491_6_g2528(.A (inc_ADD_UNS_OP5491_6_n_2636), .B
       (inc_ADD_UNS_OP5491_6_n_2633), .Q (inc_ADD_UNS_OP5491_6_n_2625));
  INX1 inc_ADD_UNS_OP5491_6_g2529(.A (inc_ADD_UNS_OP5491_6_n_2636), .Q
       (inc_ADD_UNS_OP5491_6_n_2626));
  AND4X1 inc_ADD_UNS_OP5491_6_g2530(.A (csr_minstret[30]), .B
       (csr_minstret[28]), .C (csr_minstret[31]), .D
       (csr_minstret[29]), .Q (inc_ADD_UNS_OP5491_6_n_2628));
  EO2X1 inc_ADD_UNS_OP5491_6_g2531(.A (csr_minstret[0]), .B (n_7883),
       .Q (n_7593));
  NA2X1 inc_ADD_UNS_OP5491_6_g2532(.A (csr_minstret[1]), .B
       (csr_minstret[2]), .Q (inc_ADD_UNS_OP5491_6_n_2633));
  NA2X1 inc_ADD_UNS_OP5491_6_g2533(.A (csr_minstret[0]), .B (n_7883),
       .Q (inc_ADD_UNS_OP5491_6_n_2636));
  INX1 inc_ADD_UNS_OP5491_6_g2535(.A (n_7379), .Q
       (inc_ADD_UNS_OP5491_6_n_2641));
  INX1 inc_ADD_UNS_OP5491_6_g2541(.A (n_7377), .Q
       (inc_ADD_UNS_OP5491_6_n_2657));
  OR2X2 inc_ADD_UNS_OP5491_6_g2(.A (inc_ADD_UNS_OP5491_6_n_2388), .B
       (inc_ADD_UNS_OP5491_6_n_2669), .Q (inc_ADD_UNS_OP5491_6_n_2724));
  OR2X1 inc_ADD_UNS_OP5491_6_g2556(.A (inc_ADD_UNS_OP5491_6_n_2419), .B
       (inc_ADD_UNS_OP_5_n_3760), .Q (inc_ADD_UNS_OP5491_6_n_2725));
  EO2X1 inc_ADD_UNS_OP5491_6_g2557(.A (inc_ADD_UNS_OP5491_6_n_2356), .B
       (n_7376), .Q (n_7469));
  MU2IX1 inc_ADD_UNS_OP5491_6_g2558(.S (inc_ADD_UNS_OP5491_6_n_2388),
       .IN0 (n_7381), .IN1 (inc_ADD_UNS_OP5491_6_n_2669), .Q (n_7479));
  EO2X1 inc_ADD_UNS_OP5491_6_g2559(.A (inc_ADD_UNS_OP5491_6_n_2393), .B
       (n_8571), .Q (n_7481));
  MU2IX1 inc_ADD_UNS_OP5491_6_g2560(.S (inc_ADD_UNS_OP5491_6_n_2419),
       .IN0 (n_7386), .IN1 (inc_ADD_UNS_OP_5_n_3760), .Q (n_7489));
  EO2X1 inc_ADD_UNS_OP5491_6_g2561(.A (inc_ADD_UNS_OP5491_6_n_2421), .B
       (n_7387), .Q (n_7491));
  EO2X1 inc_ADD_UNS_OP5491_6_g2562(.A (inc_ADD_UNS_OP5491_6_n_2431), .B
       (n_7389), .Q (n_7495));
  EO2X1 inc_ADD_UNS_OP5491_6_g2563(.A (inc_ADD_UNS_OP5491_6_n_2452), .B
       (n_7392), .Q (n_7501));
  EO2X1 inc_ADD_UNS_OP5491_6_g2564(.A (inc_ADD_UNS_OP5491_6_n_2468), .B
       (n_7394), .Q (n_7505));
  EN2X1 inc_ADD_UNS_OP5491_6_g2565(.A (inc_ADD_UNS_OP5491_6_n_2489), .B
       (csr_minstret[28]), .Q (n_7537));
  EN2X0 inc_ADD_UNS_OP5491_6_g2566(.A (inc_ADD_UNS_OP5491_6_n_2517), .B
       (csr_minstret[25]), .Q (n_7543));
  EN2X0 inc_ADD_UNS_OP5491_6_g2567(.A (inc_ADD_UNS_OP5491_6_n_2596), .B
       (csr_minstret[7]), .Q (n_7579));
  EN2X0 inc_ADD_UNS_OP5491_6_g2568(.A (inc_ADD_UNS_OP5491_6_n_2620), .B
       (csr_minstret[4]), .Q (n_7585));
  EO2X1 inc_ADD_UNS_OP5491_6_g2569(.A (inc_ADD_UNS_OP5491_6_n_2625), .B
       (csr_minstret[3]), .Q (n_7587));
  EN2X1 inc_ADD_UNS_OP5491_6_g2570(.A (inc_ADD_UNS_OP5491_6_n_2351), .B
       (n_7635), .Q (n_7467));
  EO2X1 inc_ADD_UNS_OP5491_6_g2571(.A (inc_ADD_UNS_OP5491_6_n_2401), .B
       (n_7384), .Q (n_7485));
  EN2X1 inc_ADD_UNS_OP5491_6_g2572(.A (inc_ADD_UNS_OP5491_6_n_2724), .B
       (n_7380), .Q (n_7477));
  EN2X1 inc_ADD_UNS_OP5491_6_g2573(.A (inc_ADD_UNS_OP5491_6_n_2446), .B
       (n_7391), .Q (n_7499));
  EO2X1 inc_ADD_UNS_OP5491_6_g2574(.A (inc_ADD_UNS_OP5491_6_n_2476), .B
       (n_7395), .Q (n_7507));
  EN2X1 inc_ADD_UNS_OP5491_6_g2575(.A (inc_ADD_UNS_OP5491_6_n_2725), .B
       (n_7385), .Q (n_7487));
  EO2X1 inc_ADD_UNS_OP5491_6_g2576(.A (inc_ADD_UNS_OP5491_6_n_2438), .B
       (n_8622), .Q (n_7497));
  EN2X1 inc_ADD_UNS_OP5491_6_g2577(.A (inc_ADD_UNS_OP5491_6_n_2440), .B
       (n_6234), .Q (n_7523));
  EO2X1 inc_ADD_UNS_OP5491_6_g2578(.A (inc_ADD_UNS_OP5491_6_n_2443), .B
       (n_6233), .Q (n_7525));
  AND6X1 inc_ADD_UNS_OP5491_6_g2580(.A (inc_ADD_UNS_OP5491_6_n_2497),
       .B (n_8354), .C (n_7395), .D (n_7394), .E (n_7398), .F (n_7397),
       .Q (inc_ADD_UNS_OP5491_6_n_2460));
  NO2I1X2 inc_ADD_UNS_OP5491_6_g2582(.B (inc_ADD_UNS_OP5491_6_n_2517),
       .AN (csr_minstret[25]), .Q (inc_ADD_UNS_OP5491_6_n_2507));
  NO2I1X2 inc_ADD_UNS_OP5491_6_g2584(.B (inc_ADD_UNS_OP5491_6_n_2489),
       .AN (csr_minstret[28]), .Q (inc_ADD_UNS_OP5491_6_n_2481));
  HAX2 inc_add_1345_58_1_g3011(.A (n_8598), .B (n_7376), .S (n_8010),
       .CO (inc_add_1345_58_1_n_3147));
  MU2IX1 inc_add_1345_58_1_g3012(.S (inc_add_1345_58_1_n_3151), .IN0
       (inc_add_1345_58_1_n_3455), .IN1 (n_7378), .Q (n_8014));
  MU2IX1 inc_add_1345_58_1_g3015(.S (inc_add_1345_58_1_n_3155), .IN0
       (inc_ADD_UNS_OP5491_6_n_2657), .IN1 (n_7377), .Q (n_8012));
  MU2IX1 inc_add_1345_58_1_g3016(.S (inc_add_1345_58_1_n_3159), .IN0
       (n_7379), .IN1 (inc_ADD_UNS_OP5491_6_n_2641), .Q (n_8016));
  NO2X1 inc_add_1345_58_1_g3017(.A (inc_add_1345_58_1_n_3159), .B
       (inc_add_1345_58_1_n_3390), .Q (inc_add_1345_58_1_n_3155));
  NO2X2 inc_add_1345_58_1_g3018(.A (inc_add_1345_58_1_n_3159), .B
       (inc_ADD_UNS_OP5491_6_n_2641), .Q (inc_add_1345_58_1_n_3151));
  NA2X2 inc_add_1345_58_1_g3021(.A (inc_add_1345_58_1_n_3166), .B
       (n_7380), .Q (inc_add_1345_58_1_n_3159));
  HAX2 inc_add_1345_58_1_g3024(.A (inc_add_1345_58_1_n_3175), .B
       (n_7381), .S (n_8020), .CO (inc_add_1345_58_1_n_3166));
  NA2X1 inc_add_1345_58_1_g3026(.A (inc_add_1345_58_1_n_3172), .B
       (n_8622), .Q (inc_add_1345_58_1_n_3169));
  HAX2 inc_add_1345_58_1_g3028(.A (inc_add_1345_58_1_n_3185), .B
       (n_7391), .S (n_8062), .CO (inc_add_1345_58_1_n_3172));
  MU2IX1 inc_add_1345_58_1_g3029(.S (inc_add_1345_58_1_n_3180), .IN0
       (n_8571), .IN1 (inc_ADD_UNS_OP_5_n_3756), .Q (n_8022));
  NO2X2 inc_add_1345_58_1_g3030(.A (inc_add_1345_58_1_n_3180), .B
       (inc_ADD_UNS_OP_5_n_3756), .Q (inc_add_1345_58_1_n_3175));
  NA2X2 inc_add_1345_58_1_g3032(.A (inc_add_1345_58_1_n_3190), .B
       (n_7383), .Q (inc_add_1345_58_1_n_3180));
  MU2IX1 inc_add_1345_58_1_g3033(.S (inc_add_1345_58_1_n_3195), .IN0
       (n_7392), .IN1 (inc_ADD_UNS_OP_5_n_3766), .Q (n_8064));
  NO2X1 inc_add_1345_58_1_g3034(.A (inc_add_1345_58_1_n_3195), .B
       (inc_ADD_UNS_OP_5_n_3766), .Q (inc_add_1345_58_1_n_3185));
  MU2IX1 inc_add_1345_58_1_g3035(.S (inc_add_1345_58_1_n_3202), .IN0
       (n_7384), .IN1 (inc_ADD_UNS_OP_5_n_3746), .Q (n_8026));
  NO2X2 inc_add_1345_58_1_g3036(.A (inc_add_1345_58_1_n_3202), .B
       (inc_ADD_UNS_OP_5_n_3746), .Q (inc_add_1345_58_1_n_3190));
  NA2X1 inc_add_1345_58_1_g3038(.A (inc_add_1345_58_1_n_3199), .B
       (n_7393), .Q (inc_add_1345_58_1_n_3195));
  HAX2 inc_add_1345_58_1_g3040(.A (inc_add_1345_58_1_n_3215), .B
       (n_7394), .S (n_8068), .CO (inc_add_1345_58_1_n_3199));
  MU2IX1 inc_add_1345_58_1_g3041(.S (inc_add_1345_58_1_n_3205), .IN0
       (inc_add_1345_58_1_n_3422), .IN1 (n_7385), .Q (n_8032));
  OR6X2 inc_add_1345_58_1_g3042(.A (inc_add_1345_58_1_n_3238), .B
       (inc_add_1345_58_1_n_3373), .C (inc_add_1345_58_1_n_3414), .D
       (n_4001), .E (n_4002), .F (inc_add_1345_58_1_n_3422), .Q
       (inc_add_1345_58_1_n_3202));
  HAX1 inc_add_1345_58_1_g3043(.A (inc_add_1345_58_1_n_3214), .B
       (n_7386), .S (n_8044), .CO (inc_add_1345_58_1_n_3205));
  NA2X1 inc_add_1345_58_1_g3045(.A (inc_add_1345_58_1_n_3210), .B
       (n_6233), .Q (inc_add_1345_58_1_n_3207));
  HAX1 inc_add_1345_58_1_g3047(.A (inc_add_1345_58_1_n_3220), .B
       (n_6235), .S (n_8092), .CO (inc_add_1345_58_1_n_3210));
  MU2IX1 inc_add_1345_58_1_g3048(.S (inc_add_1345_58_1_n_3222), .IN0
       (n_7395), .IN1 (n_8657), .Q (n_8070));
  HAX1 inc_add_1345_58_1_g3049(.A (inc_add_1345_58_1_n_3230), .B
       (n_7387), .S (n_8052), .CO (inc_add_1345_58_1_n_3214));
  NO2X1 inc_add_1345_58_1_g3050(.A (inc_add_1345_58_1_n_3222), .B
       (n_8657), .Q (inc_add_1345_58_1_n_3215));
  HAX1 inc_add_1345_58_1_g3051(.A (inc_add_1345_58_1_n_3229), .B
       (n_6236), .S (n_8094), .CO (inc_add_1345_58_1_n_3220));
  NA2X1 inc_add_1345_58_1_g3053(.A (inc_add_1345_58_1_n_3234), .B
       (n_8354), .Q (inc_add_1345_58_1_n_3222));
  EN2X1 inc_add_1345_58_1_g3055(.A (inc_add_1345_58_1_n_3236), .B
       (inc_add_1345_58_1_n_3414), .Q (n_8056));
  HAX1 inc_add_1345_58_1_g3056(.A (inc_add_1345_58_1_n_3242), .B
       (csr_mcycle[31]), .S (n_8096), .CO (inc_add_1345_58_1_n_3229));
  EN2X1 inc_add_1345_58_1_g3058(.A (inc_add_1345_58_1_n_3238), .B
       (n_7397), .Q (n_8075));
  NO2X1 inc_add_1345_58_1_g3060(.A (inc_add_1345_58_1_n_3238), .B
       (inc_add_1345_58_1_n_3373), .Q (inc_add_1345_58_1_n_3236));
  HAX2 inc_add_1345_58_1_g3063(.A (inc_add_1345_58_1_n_3248), .B
       (csr_mcycle[30]), .S (n_8098), .CO (inc_add_1345_58_1_n_3242));
  EO2X1 inc_add_1345_58_1_g3064(.A (inc_add_1345_58_1_n_3246), .B
       (n_7398), .Q (n_8077));
  OR6X2 inc_add_1345_58_1_g3065(.A (inc_add_1345_58_1_n_3267), .B
       (inc_add_1345_58_1_n_3408), .C (n_1447), .D (n_3862), .E
       (n_3863), .F (inc_add_1345_58_1_n_3434), .Q
       (inc_add_1345_58_1_n_3238));
  HAX1 inc_add_1345_58_1_g3066(.A (inc_add_1345_58_1_n_3250), .B
       (n_6238), .S (n_8080), .CO (inc_add_1345_58_1_n_3246));
  HAX2 inc_add_1345_58_1_g3067(.A (inc_add_1345_58_1_n_3252), .B
       (csr_mcycle[29]), .S (n_8100), .CO (inc_add_1345_58_1_n_3248));
  HAX1 inc_add_1345_58_1_g3068(.A (inc_add_1345_58_1_n_3254), .B
       (n_6237), .S (n_8082), .CO (inc_add_1345_58_1_n_3250));
  HAX2 inc_add_1345_58_1_g3069(.A (inc_add_1345_58_1_n_3258), .B
       (csr_mcycle[28]), .S (n_8102), .CO (inc_add_1345_58_1_n_3252));
  HAX1 inc_add_1345_58_1_g3070(.A (inc_add_1345_58_1_n_3257), .B
       (n_6232), .S (n_8084), .CO (inc_add_1345_58_1_n_3254));
  HAX1 inc_add_1345_58_1_g3072(.A (inc_add_1345_58_1_n_3266), .B
       (n_7632), .S (n_8086), .CO (inc_add_1345_58_1_n_3257));
  NO2I1X1 inc_add_1345_58_1_g3073(.B (inc_add_1345_58_1_n_3263), .AN
       (csr_mcycle[27]), .Q (inc_add_1345_58_1_n_3258));
  EO2X1 inc_add_1345_58_1_g3075(.A (inc_add_1345_58_1_n_3271), .B
       (csr_mcycle[26]), .Q (n_8106));
  NA2X1 inc_add_1345_58_1_g3076(.A (inc_add_1345_58_1_n_3271), .B
       (csr_mcycle[26]), .Q (inc_add_1345_58_1_n_3263));
  INX1 inc_add_1345_58_1_g3077(.A (inc_add_1345_58_1_n_3267), .Q
       (inc_add_1345_58_1_n_3266));
  NA5X2 inc_add_1345_58_1_g3078(.A (inc_add_1345_58_1_n_3366), .B
       (inc_add_1345_58_1_n_3280), .C (csr_mcycle[23]), .D
       (csr_mcycle[24]), .E (csr_mcycle[25]), .Q
       (inc_add_1345_58_1_n_3267));
  EO2X1 inc_add_1345_58_1_g3079(.A (inc_add_1345_58_1_n_3273), .B
       (csr_mcycle[25]), .Q (n_8108));
  HAX2 inc_add_1345_58_1_g3081(.A (inc_add_1345_58_1_n_3279), .B
       (csr_mcycle[24]), .S (n_8110), .CO (inc_add_1345_58_1_n_3273));
  EO2X1 inc_add_1345_58_1_g3082(.A (inc_add_1345_58_1_n_3280), .B
       (csr_mcycle[23]), .Q (n_8112));
  NO2I1X1 inc_add_1345_58_1_g3083(.B (inc_add_1345_58_1_n_3283), .AN
       (csr_mcycle[23]), .Q (inc_add_1345_58_1_n_3279));
  INX1 inc_add_1345_58_1_g3084(.A (inc_add_1345_58_1_n_3283), .Q
       (inc_add_1345_58_1_n_3280));
  EO2X0 inc_add_1345_58_1_g3085(.A (inc_add_1345_58_1_n_3288), .B
       (csr_mcycle[22]), .Q (n_8114));
  NA2X1 inc_add_1345_58_1_g3086(.A (inc_add_1345_58_1_n_3288), .B
       (csr_mcycle[22]), .Q (inc_add_1345_58_1_n_3283));
  EO2X0 inc_add_1345_58_1_g3087(.A (inc_add_1345_58_1_n_3293), .B
       (csr_mcycle[21]), .Q (n_8116));
  AND2X1 inc_add_1345_58_1_g3088(.A (inc_add_1345_58_1_n_3293), .B
       (csr_mcycle[21]), .Q (inc_add_1345_58_1_n_3288));
  EO2X0 inc_add_1345_58_1_g3089(.A (inc_add_1345_58_1_n_3298), .B
       (csr_mcycle[20]), .Q (n_8118));
  AND2X2 inc_add_1345_58_1_g3090(.A (inc_add_1345_58_1_n_3298), .B
       (csr_mcycle[20]), .Q (inc_add_1345_58_1_n_3293));
  EO2X1 inc_add_1345_58_1_g3091(.A (inc_add_1345_58_1_n_3301), .B
       (csr_mcycle[19]), .Q (n_8120));
  AND4X2 inc_add_1345_58_1_g3092(.A (inc_add_1345_58_1_n_3307), .B
       (csr_mcycle[17]), .C (csr_mcycle[18]), .D (csr_mcycle[19]), .Q
       (inc_add_1345_58_1_n_3298));
  HAX1 inc_add_1345_58_1_g3093(.A (inc_add_1345_58_1_n_3304), .B
       (csr_mcycle[18]), .S (n_8122), .CO (inc_add_1345_58_1_n_3301));
  HAX1 inc_add_1345_58_1_g3094(.A (inc_add_1345_58_1_n_3307), .B
       (csr_mcycle[17]), .S (n_8124), .CO (inc_add_1345_58_1_n_3304));
  HAX1 inc_add_1345_58_1_g3095(.A (inc_add_1345_58_1_n_3310), .B
       (csr_mcycle[16]), .S (n_8126), .CO (inc_add_1345_58_1_n_3307));
  NO2I1X1 inc_add_1345_58_1_g3097(.B (inc_add_1345_58_1_n_3315), .AN
       (csr_mcycle[15]), .Q (inc_add_1345_58_1_n_3310));
  EO2X1 inc_add_1345_58_1_g3099(.A (inc_add_1345_58_1_n_3320), .B
       (csr_mcycle[14]), .Q (n_8130));
  NA2X1 inc_add_1345_58_1_g3100(.A (inc_add_1345_58_1_n_3320), .B
       (csr_mcycle[14]), .Q (inc_add_1345_58_1_n_3315));
  EO2X0 inc_add_1345_58_1_g3101(.A (inc_add_1345_58_1_n_3325), .B
       (csr_mcycle[13]), .Q (n_8132));
  AND2X4 inc_add_1345_58_1_g3102(.A (inc_add_1345_58_1_n_3325), .B
       (csr_mcycle[13]), .Q (inc_add_1345_58_1_n_3320));
  NO2I1X1 inc_add_1345_58_1_g3104(.B (inc_add_1345_58_1_n_3330), .AN
       (csr_mcycle[12]), .Q (inc_add_1345_58_1_n_3325));
  EO2X0 inc_add_1345_58_1_g3106(.A (inc_add_1345_58_1_n_3335), .B
       (csr_mcycle[11]), .Q (n_8136));
  NA2X2 inc_add_1345_58_1_g3107(.A (inc_add_1345_58_1_n_3335), .B
       (csr_mcycle[11]), .Q (inc_add_1345_58_1_n_3330));
  EO2X1 inc_add_1345_58_1_g3108(.A (inc_add_1345_58_1_n_3338), .B
       (csr_mcycle[10]), .Q (n_8138));
  AND3X2 inc_add_1345_58_1_g3109(.A (inc_add_1345_58_1_n_3343), .B
       (csr_mcycle[9]), .C (csr_mcycle[10]), .Q
       (inc_add_1345_58_1_n_3335));
  HAX1 inc_add_1345_58_1_g3110(.A (inc_add_1345_58_1_n_3343), .B
       (csr_mcycle[9]), .S (n_8140), .CO (inc_add_1345_58_1_n_3338));
  NO2I1X1 inc_add_1345_58_1_g3112(.B (inc_add_1345_58_1_n_3348), .AN
       (csr_mcycle[8]), .Q (inc_add_1345_58_1_n_3343));
  EO2X0 inc_add_1345_58_1_g3114(.A (inc_add_1345_58_1_n_3353), .B
       (csr_mcycle[7]), .Q (n_8144));
  NA2X2 inc_add_1345_58_1_g3115(.A (inc_add_1345_58_1_n_3353), .B
       (csr_mcycle[7]), .Q (inc_add_1345_58_1_n_3348));
  NO2I1X2 inc_add_1345_58_1_g3117(.B (inc_add_1345_58_1_n_3358), .AN
       (csr_mcycle[6]), .Q (inc_add_1345_58_1_n_3353));
  EO2X0 inc_add_1345_58_1_g3119(.A (inc_add_1345_58_1_n_3370), .B
       (csr_mcycle[5]), .Q (n_8148));
  NA2X2 inc_add_1345_58_1_g3120(.A (inc_add_1345_58_1_n_3370), .B
       (csr_mcycle[5]), .Q (inc_add_1345_58_1_n_3358));
  EO2X1 inc_add_1345_58_1_g3121(.A (inc_add_1345_58_1_n_3364), .B
       (csr_mcycle[3]), .Q (n_8152));
  HAX1 inc_add_1345_58_1_g3122(.A (inc_add_1345_58_1_n_3399), .B
       (csr_mcycle[2]), .S (n_8154), .CO (inc_add_1345_58_1_n_3364));
  EN2X0 inc_add_1345_58_1_g3123(.A (n_8597), .B (csr_mcycle[4]), .Q
       (n_8150));
  AND5X1 inc_add_1345_58_1_g3124(.A (n_6233), .B (n_6234), .C (n_6236),
       .D (n_6235), .E (inc_add_1345_58_1_n_3382), .Q
       (inc_add_1345_58_1_n_3366));
  NO2I1X2 inc_add_1345_58_1_g3125(.B (n_8597), .AN (csr_mcycle[4]), .Q
       (inc_add_1345_58_1_n_3370));
  NA3X1 inc_add_1345_58_1_g3126(.A (inc_add_1345_58_1_n_3378), .B
       (inc_add_1345_58_1_n_3387), .C (n_7392), .Q
       (inc_add_1345_58_1_n_3373));
  AND5X1 inc_add_1345_58_1_g3128(.A (n_7391), .B (n_8354), .C (n_7394),
       .D (n_7393), .E (n_7395), .Q (inc_add_1345_58_1_n_3378));
  AND6X1 inc_add_1345_58_1_g3129(.A (csr_mcycle[26]), .B
       (csr_mcycle[30]), .C (csr_mcycle[27]), .D (csr_mcycle[29]), .E
       (csr_mcycle[28]), .F (csr_mcycle[31]), .Q
       (inc_add_1345_58_1_n_3382));
  AND3X1 inc_add_1345_58_1_g3130(.A (n_8622), .B (n_7397), .C (n_7389),
       .Q (inc_add_1345_58_1_n_3387));
  EO2X1 inc_add_1345_58_1_g3131(.A (csr_mcycle[0]), .B (csr_mcycle[1]),
       .Q (n_8156));
  NA2X1 inc_add_1345_58_1_g3132(.A (n_7379), .B (n_7378), .Q
       (inc_add_1345_58_1_n_3390));
  AND2X1 inc_add_1345_58_1_g3135(.A (csr_mcycle[0]), .B
       (csr_mcycle[1]), .Q (inc_add_1345_58_1_n_3399));
  INX1 inc_add_1345_58_1_g3139(.A (n_6237), .Q
       (inc_add_1345_58_1_n_3408));
  INX1 inc_add_1345_58_1_g3142(.A (n_7388), .Q
       (inc_add_1345_58_1_n_3414));
  INX1 inc_add_1345_58_1_g3146(.A (n_7385), .Q
       (inc_add_1345_58_1_n_3422));
  INX1 inc_add_1345_58_1_g3152(.A (n_6232), .Q
       (inc_add_1345_58_1_n_3434));
  EO2X1 inc_add_1345_58_1_g2(.A (inc_add_1345_58_1_n_3166), .B
       (n_7380), .Q (n_8018));
  EO2X1 inc_add_1345_58_1_g3160(.A (inc_add_1345_58_1_n_3172), .B
       (n_8622), .Q (n_8060));
  EO2X1 inc_add_1345_58_1_g3161(.A (inc_add_1345_58_1_n_3210), .B
       (n_6233), .Q (n_8090));
  EO2X1 inc_add_1345_58_1_g3162(.A (inc_add_1345_58_1_n_3234), .B
       (n_8354), .Q (n_8072));
  EN2X1 inc_add_1345_58_1_g3163(.A (inc_add_1345_58_1_n_3263), .B
       (csr_mcycle[27]), .Q (n_8104));
  EN2X0 inc_add_1345_58_1_g3164(.A (inc_add_1345_58_1_n_3315), .B
       (csr_mcycle[15]), .Q (n_8128));
  EN2X0 inc_add_1345_58_1_g3165(.A (inc_add_1345_58_1_n_3330), .B
       (csr_mcycle[12]), .Q (n_8134));
  EN2X0 inc_add_1345_58_1_g3166(.A (inc_add_1345_58_1_n_3348), .B
       (csr_mcycle[8]), .Q (n_8142));
  EN2X0 inc_add_1345_58_1_g3167(.A (inc_add_1345_58_1_n_3358), .B
       (csr_mcycle[6]), .Q (n_8146));
  EO2X1 inc_add_1345_58_1_g3168(.A (inc_add_1345_58_1_n_3147), .B
       (n_7635), .Q (n_8008));
  EO2X1 inc_add_1345_58_1_g3169(.A (inc_add_1345_58_1_n_3190), .B
       (n_7383), .Q (n_8024));
  EN2X1 inc_add_1345_58_1_g3170(.A (inc_add_1345_58_1_n_3207), .B
       (n_6234), .Q (n_8088));
  EN2X1 inc_add_1345_58_1_g3171(.A (inc_add_1345_58_1_n_3169), .B
       (n_7389), .Q (n_8058));
  EO2X1 inc_add_1345_58_1_g3172(.A (inc_add_1345_58_1_n_3199), .B
       (n_7393), .Q (n_8066));
  AND2X1 inc_add_1345_58_1_g3176(.A (inc_add_1345_58_1_n_3236), .B
       (n_7388), .Q (inc_add_1345_58_1_n_3230));
  NO2I1X1 inc_add_1345_58_1_g3178(.B (inc_add_1345_58_1_n_3238), .AN
       (n_7397), .Q (inc_add_1345_58_1_n_3234));
  AND2X1 inc_add_1345_58_1_g3182(.A (inc_add_1345_58_1_n_3273), .B
       (csr_mcycle[25]), .Q (inc_add_1345_58_1_n_3271));
  NA2X2 inc_add_1347_34_2_g2343(.A (inc_add_1347_34_2_n_2321), .B
       (csr_mcycle[62]), .Q (inc_add_1347_34_2_n_2311));
  NA2X2 inc_add_1347_34_2_g2346(.A (inc_add_1347_34_2_n_2326), .B
       (csr_mcycle[54]), .Q (inc_add_1347_34_2_n_2316));
  MU2IX1 inc_add_1347_34_2_g2348(.S (inc_add_1347_34_2_n_2331), .IN0
       (csr_mcycle[61]), .IN1 (inc_add_1347_34_2_n_2589), .Q (n_8011));
  NO2X2 inc_add_1347_34_2_g2349(.A (inc_add_1347_34_2_n_2331), .B
       (inc_add_1347_34_2_n_2589), .Q (inc_add_1347_34_2_n_2321));
  MU2IX1 inc_add_1347_34_2_g2350(.S (inc_add_1347_34_2_n_2336), .IN0
       (csr_mcycle[53]), .IN1 (inc_add_1347_34_2_n_2595), .Q (n_8027));
  NO2X4 inc_add_1347_34_2_g2351(.A (inc_add_1347_34_2_n_2336), .B
       (inc_add_1347_34_2_n_2595), .Q (inc_add_1347_34_2_n_2326));
  NA2X2 inc_add_1347_34_2_g2353(.A (inc_add_1347_34_2_n_2341), .B
       (csr_mcycle[60]), .Q (inc_add_1347_34_2_n_2331));
  NA2X1 inc_add_1347_34_2_g2356(.A (inc_add_1347_34_2_n_2347), .B
       (csr_mcycle[52]), .Q (inc_add_1347_34_2_n_2336));
  MU2IX1 inc_add_1347_34_2_g2358(.S (inc_add_1347_34_2_n_2352), .IN0
       (csr_mcycle[59]), .IN1 (inc_add_1343_59_4_n_3758), .Q (n_8015));
  NO2X2 inc_add_1347_34_2_g2360(.A (inc_add_1347_34_2_n_2352), .B
       (inc_add_1343_59_4_n_3758), .Q (inc_add_1347_34_2_n_2341));
  MU2IX1 inc_add_1347_34_2_g2361(.S (inc_add_1347_34_2_n_2357), .IN0
       (csr_mcycle[51]), .IN1 (inc_add_1343_59_4_n_3788), .Q (n_8050));
  NO2X4 inc_add_1347_34_2_g2362(.A (inc_add_1347_34_2_n_2357), .B
       (inc_add_1343_59_4_n_3788), .Q (inc_add_1347_34_2_n_2347));
  NA2X1 inc_add_1347_34_2_g2364(.A (inc_add_1347_34_2_n_2362), .B
       (csr_mcycle[58]), .Q (inc_add_1347_34_2_n_2352));
  NA2X2 inc_add_1347_34_2_g2367(.A (inc_add_1347_34_2_n_2368), .B
       (csr_mcycle[50]), .Q (inc_add_1347_34_2_n_2357));
  MU2IX1 inc_add_1347_34_2_g2369(.S (inc_add_1347_34_2_n_2373), .IN0
       (csr_mcycle[57]), .IN1 (inc_add_1343_59_4_n_3775), .Q (n_8019));
  NO2X2 inc_add_1347_34_2_g2371(.A (inc_add_1347_34_2_n_2373), .B
       (inc_add_1343_59_4_n_3775), .Q (inc_add_1347_34_2_n_2362));
  MU2IX1 inc_add_1347_34_2_g2372(.S (inc_add_1347_34_2_n_2650), .IN0
       (csr_mcycle[49]), .IN1 (inc_add_1343_59_4_n_3784), .Q (n_8057));
  NO2X2 inc_add_1347_34_2_g2373(.A (inc_add_1347_34_2_n_2650), .B
       (inc_add_1343_59_4_n_3784), .Q (inc_add_1347_34_2_n_2368));
  NA2X2 inc_add_1347_34_2_g2375(.A (inc_add_1347_34_2_n_2377), .B
       (csr_mcycle[56]), .Q (inc_add_1347_34_2_n_2373));
  NO2X2 inc_add_1347_34_2_g2378(.A (inc_add_1347_34_2_n_2381), .B
       (inc_add_1347_34_2_n_2544), .Q (inc_add_1347_34_2_n_2377));
  NA6X2 inc_add_1347_34_2_g2383(.A (inc_add_1347_34_2_n_2401), .B
       (csr_mcycle[43]), .C (csr_mcycle[45]), .D (csr_mcycle[44]), .E
       (csr_mcycle[46]), .F (csr_mcycle[47]), .Q
       (inc_add_1347_34_2_n_2381));
  NA2X1 inc_add_1347_34_2_g2385(.A (inc_add_1347_34_2_n_2391), .B
       (csr_mcycle[46]), .Q (inc_add_1347_34_2_n_2389));
  HAX2 inc_add_1347_34_2_g2387(.A (inc_add_1347_34_2_n_2396), .B
       (csr_mcycle[45]), .S (n_8065), .CO (inc_add_1347_34_2_n_2391));
  EN2X1 inc_add_1347_34_2_g2388(.A (inc_add_1347_34_2_n_2400), .B
       (csr_mcycle[44]), .Q (n_8067));
  EO2X1 inc_add_1347_34_2_g2390(.A (inc_add_1347_34_2_n_2401), .B
       (csr_mcycle[43]), .Q (n_8069));
  NA2X1 inc_add_1347_34_2_g2391(.A (inc_add_1347_34_2_n_2401), .B
       (csr_mcycle[43]), .Q (inc_add_1347_34_2_n_2400));
  EO2X1 inc_add_1347_34_2_g2393(.A (inc_add_1347_34_2_n_2409), .B
       (csr_mcycle[42]), .Q (n_8071));
  AND6X2 inc_add_1347_34_2_g2394(.A (inc_add_1347_34_2_n_2422), .B
       (csr_mcycle[38]), .C (csr_mcycle[40]), .D (csr_mcycle[39]), .E
       (csr_mcycle[41]), .F (csr_mcycle[42]), .Q
       (inc_add_1347_34_2_n_2401));
  HAX1 inc_add_1347_34_2_g2395(.A (inc_add_1347_34_2_n_2411), .B
       (csr_mcycle[41]), .S (n_8074), .CO (inc_add_1347_34_2_n_2409));
  HAX1 inc_add_1347_34_2_g2396(.A (inc_add_1347_34_2_n_2413), .B
       (csr_mcycle[40]), .S (n_8076), .CO (inc_add_1347_34_2_n_2411));
  HAX2 inc_add_1347_34_2_g2397(.A (inc_add_1347_34_2_n_2417), .B
       (csr_mcycle[39]), .S (n_8079), .CO (inc_add_1347_34_2_n_2413));
  HAX2 inc_add_1347_34_2_g2398(.A (inc_add_1347_34_2_n_2422), .B
       (csr_mcycle[38]), .S (n_8081), .CO (inc_add_1347_34_2_n_2417));
  EO2X1 inc_add_1347_34_2_g2399(.A (inc_add_1347_34_2_n_2426), .B
       (csr_mcycle[37]), .Q (n_8083));
  AND6X2 inc_add_1347_34_2_g2400(.A (inc_add_1347_34_2_n_2446), .B
       (csr_mcycle[33]), .C (csr_mcycle[35]), .D (csr_mcycle[34]), .E
       (csr_mcycle[36]), .F (csr_mcycle[37]), .Q
       (inc_add_1347_34_2_n_2422));
  EO2X1 inc_add_1347_34_2_g2401(.A (inc_add_1347_34_2_n_2429), .B
       (csr_mcycle[28]), .Q (n_8101));
  HAX1 inc_add_1347_34_2_g2402(.A (inc_add_1347_34_2_n_2431), .B
       (csr_mcycle[36]), .S (n_8085), .CO (inc_add_1347_34_2_n_2426));
  HAX1 inc_add_1347_34_2_g2403(.A (inc_add_1347_34_2_n_2434), .B
       (csr_mcycle[27]), .S (n_8103), .CO (inc_add_1347_34_2_n_2429));
  HAX1 inc_add_1347_34_2_g2404(.A (inc_add_1347_34_2_n_2436), .B
       (csr_mcycle[35]), .S (n_8087), .CO (inc_add_1347_34_2_n_2431));
  HAX1 inc_add_1347_34_2_g2405(.A (inc_add_1347_34_2_n_2439), .B
       (csr_mcycle[26]), .S (n_8105), .CO (inc_add_1347_34_2_n_2434));
  HAX1 inc_add_1347_34_2_g2406(.A (inc_add_1347_34_2_n_2441), .B
       (csr_mcycle[34]), .S (n_8089), .CO (inc_add_1347_34_2_n_2436));
  HAX1 inc_add_1347_34_2_g2407(.A (inc_add_1347_34_2_n_2445), .B
       (csr_mcycle[25]), .S (n_8107), .CO (inc_add_1347_34_2_n_2439));
  HAX1 inc_add_1347_34_2_g2408(.A (inc_add_1347_34_2_n_2446), .B
       (csr_mcycle[33]), .S (n_8091), .CO (inc_add_1347_34_2_n_2441));
  HAX1 inc_add_1347_34_2_g2409(.A (inc_add_1347_34_2_n_2449), .B
       (csr_mcycle[24]), .S (n_8109), .CO (inc_add_1347_34_2_n_2445));
  HAX2 inc_add_1347_34_2_g2410(.A (inc_add_1347_34_2_n_2451), .B
       (csr_mcycle[32]), .S (n_8093), .CO (inc_add_1347_34_2_n_2446));
  HAX1 inc_add_1347_34_2_g2411(.A (inc_add_1347_34_2_n_2453), .B
       (csr_mcycle[23]), .S (n_8111), .CO (inc_add_1347_34_2_n_2449));
  HAX2 inc_add_1347_34_2_g2412(.A (inc_add_1347_34_2_n_2455), .B
       (csr_mcycle[31]), .S (n_8095), .CO (inc_add_1347_34_2_n_2451));
  HAX1 inc_add_1347_34_2_g2413(.A (inc_add_1347_34_2_n_2457), .B
       (csr_mcycle[22]), .S (n_8113), .CO (inc_add_1347_34_2_n_2453));
  HAX2 inc_add_1347_34_2_g2414(.A (inc_add_1347_34_2_n_2459), .B
       (csr_mcycle[30]), .S (n_8097), .CO (inc_add_1347_34_2_n_2455));
  HAX1 inc_add_1347_34_2_g2415(.A (inc_add_1347_34_2_n_2461), .B
       (csr_mcycle[21]), .S (n_8115), .CO (inc_add_1347_34_2_n_2457));
  HAX2 inc_add_1347_34_2_g2416(.A (inc_add_1347_34_2_n_2462), .B
       (csr_mcycle[29]), .S (n_8099), .CO (inc_add_1347_34_2_n_2459));
  HAX1 inc_add_1347_34_2_g2417(.A (inc_add_1347_34_2_n_2464), .B
       (csr_mcycle[20]), .S (n_8117), .CO (inc_add_1347_34_2_n_2461));
  AND5X1 inc_add_1347_34_2_g2418(.A (inc_add_1347_34_2_n_2472), .B
       (inc_add_1347_34_2_n_2547), .C (inc_add_1347_34_2_n_2553), .D
       (csr_mcycle[18]), .E (csr_mcycle[19]), .Q
       (inc_add_1347_34_2_n_2462));
  HAX1 inc_add_1347_34_2_g2419(.A (inc_add_1347_34_2_n_2467), .B
       (csr_mcycle[19]), .S (n_8119), .CO (inc_add_1347_34_2_n_2464));
  HAX1 inc_add_1347_34_2_g2420(.A (inc_add_1347_34_2_n_2472), .B
       (csr_mcycle[18]), .S (n_8121), .CO (inc_add_1347_34_2_n_2467));
  EO2X0 inc_add_1347_34_2_g2421(.A (inc_add_1347_34_2_n_2652), .B
       (csr_mcycle[17]), .Q (n_8123));
  AND2X4 inc_add_1347_34_2_g2422(.A (inc_add_1347_34_2_n_2652), .B
       (csr_mcycle[17]), .Q (inc_add_1347_34_2_n_2472));
  EO2X0 inc_add_1347_34_2_g2423(.A (inc_add_1347_34_2_n_2482), .B
       (csr_mcycle[16]), .Q (n_8125));
  NO2I1X2 inc_add_1347_34_2_g2427(.B (inc_add_1347_34_2_n_2487), .AN
       (csr_mcycle[15]), .Q (inc_add_1347_34_2_n_2482));
  EO2X0 inc_add_1347_34_2_g2429(.A (inc_add_1347_34_2_n_2492), .B
       (csr_mcycle[14]), .Q (n_8129));
  NA2X2 inc_add_1347_34_2_g2430(.A (inc_add_1347_34_2_n_2492), .B
       (csr_mcycle[14]), .Q (inc_add_1347_34_2_n_2487));
  NO2I1X1 inc_add_1347_34_2_g2432(.B (inc_add_1347_34_2_n_2497), .AN
       (csr_mcycle[13]), .Q (inc_add_1347_34_2_n_2492));
  EO2X0 inc_add_1347_34_2_g2434(.A (inc_add_1347_34_2_n_2502), .B
       (csr_mcycle[12]), .Q (n_8133));
  NA2X2 inc_add_1347_34_2_g2435(.A (inc_add_1347_34_2_n_2502), .B
       (csr_mcycle[12]), .Q (inc_add_1347_34_2_n_2497));
  EO2X1 inc_add_1347_34_2_g2436(.A (inc_add_1347_34_2_n_2505), .B
       (csr_mcycle[11]), .Q (n_8135));
  AND3X2 inc_add_1347_34_2_g2437(.A (inc_add_1347_34_2_n_2510), .B
       (csr_mcycle[10]), .C (csr_mcycle[11]), .Q
       (inc_add_1347_34_2_n_2502));
  HAX1 inc_add_1347_34_2_g2438(.A (inc_add_1347_34_2_n_2510), .B
       (csr_mcycle[10]), .S (n_8137), .CO (inc_add_1347_34_2_n_2505));
  EO2X0 inc_add_1347_34_2_g2439(.A (inc_add_1347_34_2_n_2515), .B
       (csr_mcycle[9]), .Q (n_8139));
  AND2X2 inc_add_1347_34_2_g2440(.A (inc_add_1347_34_2_n_2515), .B
       (csr_mcycle[9]), .Q (inc_add_1347_34_2_n_2510));
  NO2I1X1 inc_add_1347_34_2_g2442(.B (inc_add_1347_34_2_n_2520), .AN
       (csr_mcycle[8]), .Q (inc_add_1347_34_2_n_2515));
  EO2X0 inc_add_1347_34_2_g2444(.A (inc_add_1347_34_2_n_2525), .B
       (csr_mcycle[7]), .Q (n_8143));
  NA2X2 inc_add_1347_34_2_g2445(.A (inc_add_1347_34_2_n_2525), .B
       (csr_mcycle[7]), .Q (inc_add_1347_34_2_n_2520));
  NO2I1X2 inc_add_1347_34_2_g2447(.B (inc_add_1347_34_2_n_2530), .AN
       (csr_mcycle[6]), .Q (inc_add_1347_34_2_n_2525));
  EO2X0 inc_add_1347_34_2_g2449(.A (inc_add_1347_34_2_n_2538), .B
       (csr_mcycle[5]), .Q (n_8147));
  NA2X2 inc_add_1347_34_2_g2450(.A (inc_add_1347_34_2_n_2538), .B
       (csr_mcycle[5]), .Q (inc_add_1347_34_2_n_2530));
  EO2X1 inc_add_1347_34_2_g2451(.A (inc_add_1347_34_2_n_2536), .B
       (csr_mcycle[3]), .Q (n_8151));
  HAX1 inc_add_1347_34_2_g2452(.A (inc_add_1347_34_2_n_2561), .B
       (csr_mcycle[2]), .S (n_8153), .CO (inc_add_1347_34_2_n_2536));
  EN2X0 inc_add_1347_34_2_g2453(.A (n_8599), .B (csr_mcycle[4]), .Q
       (n_8149));
  NO2I1X2 inc_add_1347_34_2_g2454(.B (n_8599), .AN (csr_mcycle[4]), .Q
       (inc_add_1347_34_2_n_2538));
  NA5X1 inc_add_1347_34_2_g2456(.A (inc_add_1347_34_2_n_2558), .B
       (csr_mcycle[48]), .C (csr_mcycle[49]), .D (csr_mcycle[53]), .E
       (csr_mcycle[52]), .Q (inc_add_1347_34_2_n_2544));
  AND5X1 inc_add_1347_34_2_g2457(.A (csr_mcycle[27]), .B
       (csr_mcycle[28]), .C (csr_mcycle[21]), .D (csr_mcycle[20]), .E
       (csr_mcycle[22]), .Q (inc_add_1347_34_2_n_2547));
  AND4X1 inc_add_1347_34_2_g2458(.A (csr_mcycle[25]), .B
       (csr_mcycle[23]), .C (csr_mcycle[26]), .D (csr_mcycle[24]), .Q
       (inc_add_1347_34_2_n_2553));
  AND4X1 inc_add_1347_34_2_g2459(.A (csr_mcycle[54]), .B
       (csr_mcycle[50]), .C (csr_mcycle[55]), .D (csr_mcycle[51]), .Q
       (inc_add_1347_34_2_n_2558));
  EO2X0 inc_add_1347_34_2_g2460(.A (csr_mcycle[0]), .B (csr_mcycle[1]),
       .Q (n_8155));
  AND2X1 inc_add_1347_34_2_g2461(.A (csr_mcycle[0]), .B
       (csr_mcycle[1]), .Q (inc_add_1347_34_2_n_2561));
  INX1 inc_add_1347_34_2_g2465(.A (csr_mcycle[61]), .Q
       (inc_add_1347_34_2_n_2589));
  INX1 inc_add_1347_34_2_g2467(.A (csr_mcycle[53]), .Q
       (inc_add_1347_34_2_n_2595));
  EO2X1 inc_add_1347_34_2_g2(.A (inc_add_1347_34_2_n_2321), .B
       (csr_mcycle[62]), .Q (n_8009));
  EO2X1 inc_add_1347_34_2_g2479(.A (inc_add_1347_34_2_n_2326), .B
       (csr_mcycle[54]), .Q (n_8025));
  EO2X1 inc_add_1347_34_2_g2480(.A (inc_add_1347_34_2_n_2341), .B
       (csr_mcycle[60]), .Q (n_8013));
  EO2X1 inc_add_1347_34_2_g2481(.A (inc_add_1347_34_2_n_2347), .B
       (csr_mcycle[52]), .Q (n_8038));
  EO2X1 inc_add_1347_34_2_g2482(.A (inc_add_1347_34_2_n_2362), .B
       (csr_mcycle[58]), .Q (n_8017));
  EO2X1 inc_add_1347_34_2_g2483(.A (inc_add_1347_34_2_n_2368), .B
       (csr_mcycle[50]), .Q (n_8055));
  EO2X1 inc_add_1347_34_2_g2484(.A (inc_add_1347_34_2_n_2377), .B
       (csr_mcycle[56]), .Q (n_8021));
  NA2I1X1 inc_add_1347_34_2_g2485(.B (csr_mcycle[48]), .AN
       (inc_add_1347_34_2_n_2381), .Q (inc_add_1347_34_2_n_2650));
  EO2X1 inc_add_1347_34_2_g2486(.A (inc_add_1347_34_2_n_2391), .B
       (csr_mcycle[46]), .Q (n_8063));
  AND2X1 inc_add_1347_34_2_g2487(.A (inc_add_1347_34_2_n_2482), .B
       (csr_mcycle[16]), .Q (inc_add_1347_34_2_n_2652));
  EN2X0 inc_add_1347_34_2_g2488(.A (inc_add_1347_34_2_n_2487), .B
       (csr_mcycle[15]), .Q (n_8127));
  EN2X0 inc_add_1347_34_2_g2489(.A (inc_add_1347_34_2_n_2497), .B
       (csr_mcycle[13]), .Q (n_8131));
  EN2X0 inc_add_1347_34_2_g2490(.A (inc_add_1347_34_2_n_2520), .B
       (csr_mcycle[8]), .Q (n_8141));
  EN2X0 inc_add_1347_34_2_g2491(.A (inc_add_1347_34_2_n_2530), .B
       (csr_mcycle[6]), .Q (n_8145));
  EN2X1 inc_add_1347_34_2_g2492(.A (inc_add_1347_34_2_n_2389), .B
       (csr_mcycle[47]), .Q (n_8061));
  EN2X1 inc_add_1347_34_2_g2493(.A (inc_add_1347_34_2_n_2381), .B
       (csr_mcycle[48]), .Q (n_8059));
  AND6X1 inc_add_1347_34_2_g2497(.A (inc_add_1347_34_2_n_2413), .B
       (csr_mcycle[40]), .C (csr_mcycle[42]), .D (csr_mcycle[41]), .E
       (csr_mcycle[43]), .F (csr_mcycle[44]), .Q
       (inc_add_1347_34_2_n_2396));
  NA2X2 inc_ADD_UNS_OP5492_3_g2371(.A (inc_ADD_UNS_OP5492_3_n_2339), .B
       (csr_minstret[62]), .Q (inc_ADD_UNS_OP5492_3_n_2334));
  MU2IX1 inc_ADD_UNS_OP5492_3_g2373(.S (inc_ADD_UNS_OP5492_3_n_2344),
       .IN0 (csr_minstret[61]), .IN1 (inc_ADD_UNS_OP5492_3_n_2647), .Q
       (n_7470));
  NO2X4 inc_ADD_UNS_OP5492_3_g2374(.A (inc_ADD_UNS_OP5492_3_n_2344), .B
       (inc_ADD_UNS_OP5492_3_n_2647), .Q (inc_ADD_UNS_OP5492_3_n_2339));
  NA2X4 inc_ADD_UNS_OP5492_3_g2376(.A (inc_ADD_UNS_OP5492_3_n_2350), .B
       (csr_minstret[60]), .Q (inc_ADD_UNS_OP5492_3_n_2344));
  MU2IX1 inc_ADD_UNS_OP5492_3_g2379(.S (inc_ADD_UNS_OP5492_3_n_2361),
       .IN0 (csr_minstret[59]), .IN1 (inc_ADD_UNS_OP5492_3_n_2649), .Q
       (n_7474));
  NO2X4 inc_ADD_UNS_OP5492_3_g2381(.A (inc_ADD_UNS_OP5492_3_n_2361), .B
       (inc_ADD_UNS_OP5492_3_n_2649), .Q (inc_ADD_UNS_OP5492_3_n_2350));
  NA2X1 inc_ADD_UNS_OP5492_3_g2383(.A (inc_ADD_UNS_OP5492_3_n_2366), .B
       (csr_minstret[51]), .Q (inc_ADD_UNS_OP5492_3_n_2356));
  NA2X2 inc_ADD_UNS_OP5492_3_g2386(.A (inc_ADD_UNS_OP5492_3_n_2371), .B
       (csr_minstret[58]), .Q (inc_ADD_UNS_OP5492_3_n_2361));
  MU2IX1 inc_ADD_UNS_OP5492_3_g2387(.S (inc_ADD_UNS_OP5492_3_n_2377),
       .IN0 (csr_minstret[50]), .IN1 (inc_ADD_UNS_OP5492_3_n_2615), .Q
       (n_7492));
  NO2X2 inc_ADD_UNS_OP5492_3_g2389(.A (inc_ADD_UNS_OP5492_3_n_2377), .B
       (inc_ADD_UNS_OP5492_3_n_2615), .Q (inc_ADD_UNS_OP5492_3_n_2366));
  MU2IX1 inc_ADD_UNS_OP5492_3_g2390(.S (inc_ADD_UNS_OP5492_3_n_2383),
       .IN0 (csr_minstret[57]), .IN1 (inc_ADD_UNS_OP5492_3_n_2656), .Q
       (n_7478));
  NO2X4 inc_ADD_UNS_OP5492_3_g2392(.A (inc_ADD_UNS_OP5492_3_n_2383), .B
       (inc_ADD_UNS_OP5492_3_n_2656), .Q (inc_ADD_UNS_OP5492_3_n_2371));
  NA2X2 inc_ADD_UNS_OP5492_3_g2394(.A (inc_ADD_UNS_OP5492_3_n_2380), .B
       (csr_minstret[49]), .Q (inc_ADD_UNS_OP5492_3_n_2377));
  HAX2 inc_ADD_UNS_OP5492_3_g2396(.A (inc_ADD_UNS_OP5492_3_n_2394), .B
       (csr_minstret[48]), .S (n_7496), .CO
       (inc_ADD_UNS_OP5492_3_n_2380));
  NA2X4 inc_ADD_UNS_OP5492_3_g2398(.A (inc_ADD_UNS_OP5492_3_n_2388), .B
       (csr_minstret[56]), .Q (inc_ADD_UNS_OP5492_3_n_2383));
  MU2IX1 inc_ADD_UNS_OP5492_3_g2400(.S (inc_ADD_UNS_OP5492_3_n_2399),
       .IN0 (csr_minstret[55]), .IN1 (inc_ADD_UNS_OP5492_3_n_2608), .Q
       (n_7482));
  NO2X2 inc_ADD_UNS_OP5492_3_g2402(.A (inc_ADD_UNS_OP5492_3_n_2399), .B
       (inc_ADD_UNS_OP5492_3_n_2608), .Q (inc_ADD_UNS_OP5492_3_n_2388));
  MU2IX1 inc_ADD_UNS_OP5492_3_g2403(.S (inc_ADD_UNS_OP5492_3_n_2404),
       .IN0 (csr_minstret[47]), .IN1 (inc_ADD_UNS_OP_5_n_3838), .Q
       (n_7498));
  NO2X2 inc_ADD_UNS_OP5492_3_g2404(.A (inc_ADD_UNS_OP5492_3_n_2404), .B
       (inc_ADD_UNS_OP_5_n_3838), .Q (inc_ADD_UNS_OP5492_3_n_2394));
  NA2X2 inc_ADD_UNS_OP5492_3_g2406(.A (inc_ADD_UNS_OP5492_3_n_2409), .B
       (csr_minstret[54]), .Q (inc_ADD_UNS_OP5492_3_n_2399));
  NA2X1 inc_ADD_UNS_OP5492_3_g2409(.A (inc_ADD_UNS_OP5492_3_n_2413), .B
       (csr_minstret[46]), .Q (inc_ADD_UNS_OP5492_3_n_2404));
  AND6X2 inc_ADD_UNS_OP5492_3_g2413(.A (inc_ADD_UNS_OP5492_3_n_2431),
       .B (inc_ADD_UNS_OP5492_3_n_2571), .C (csr_minstret[42]), .D
       (csr_minstret[44]), .E (csr_minstret[43]), .F
       (csr_minstret[53]), .Q (inc_ADD_UNS_OP5492_3_n_2409));
  MU2IX1 inc_ADD_UNS_OP5492_3_g2414(.S (inc_ADD_UNS_OP5492_3_n_2419),
       .IN0 (csr_minstret[45]), .IN1 (inc_ADD_UNS_OP5492_3_n_2613), .Q
       (n_7502));
  NO2X2 inc_ADD_UNS_OP5492_3_g2415(.A (inc_ADD_UNS_OP5492_3_n_2419), .B
       (inc_ADD_UNS_OP5492_3_n_2613), .Q (inc_ADD_UNS_OP5492_3_n_2413));
  NA6X2 inc_ADD_UNS_OP5492_3_g2420(.A (inc_ADD_UNS_OP5492_3_n_2444), .B
       (csr_minstret[40]), .C (csr_minstret[42]), .D
       (csr_minstret[41]), .E (csr_minstret[43]), .F
       (csr_minstret[44]), .Q (inc_ADD_UNS_OP5492_3_n_2419));
  NA3X1 inc_ADD_UNS_OP5492_3_g2422(.A (inc_ADD_UNS_OP5492_3_n_2431), .B
       (csr_minstret[42]), .C (csr_minstret[43]), .Q
       (inc_ADD_UNS_OP5492_3_n_2427));
  EO2X1 inc_ADD_UNS_OP5492_3_g2423(.A (inc_ADD_UNS_OP5492_3_n_2431), .B
       (csr_minstret[42]), .Q (n_7508));
  NA2X1 inc_ADD_UNS_OP5492_3_g2424(.A (inc_ADD_UNS_OP5492_3_n_2431), .B
       (csr_minstret[42]), .Q (inc_ADD_UNS_OP5492_3_n_2430));
  AND6X2 inc_ADD_UNS_OP5492_3_g2428(.A (inc_ADD_UNS_OP5492_3_n_2455),
       .B (csr_minstret[37]), .C (csr_minstret[39]), .D
       (csr_minstret[38]), .E (csr_minstret[40]), .F
       (csr_minstret[41]), .Q (inc_ADD_UNS_OP5492_3_n_2431));
  HAX1 inc_ADD_UNS_OP5492_3_g2429(.A (inc_ADD_UNS_OP5492_3_n_2444), .B
       (csr_minstret[40]), .S (n_7512), .CO
       (inc_ADD_UNS_OP5492_3_n_2439));
  EO2X1 inc_ADD_UNS_OP5492_3_g2430(.A (inc_ADD_UNS_OP5492_3_n_2448), .B
       (csr_minstret[39]), .Q (n_7514));
  AND6X2 inc_ADD_UNS_OP5492_3_g2431(.A (inc_ADD_UNS_OP5492_3_n_2468),
       .B (csr_minstret[35]), .C (csr_minstret[37]), .D
       (csr_minstret[36]), .E (csr_minstret[38]), .F
       (csr_minstret[39]), .Q (inc_ADD_UNS_OP5492_3_n_2444));
  HAX1 inc_ADD_UNS_OP5492_3_g2432(.A (inc_ADD_UNS_OP5492_3_n_2450), .B
       (csr_minstret[38]), .S (n_7516), .CO
       (inc_ADD_UNS_OP5492_3_n_2448));
  HAX1 inc_ADD_UNS_OP5492_3_g2433(.A (inc_ADD_UNS_OP5492_3_n_2455), .B
       (csr_minstret[37]), .S (n_7518), .CO
       (inc_ADD_UNS_OP5492_3_n_2450));
  EO2X1 inc_ADD_UNS_OP5492_3_g2434(.A (inc_ADD_UNS_OP5492_3_n_2459), .B
       (csr_minstret[36]), .Q (n_7520));
  AND6X2 inc_ADD_UNS_OP5492_3_g2435(.A (inc_ADD_UNS_OP5492_3_n_2480),
       .B (csr_minstret[32]), .C (csr_minstret[34]), .D
       (csr_minstret[33]), .E (csr_minstret[35]), .F
       (csr_minstret[36]), .Q (inc_ADD_UNS_OP5492_3_n_2455));
  EO2X1 inc_ADD_UNS_OP5492_3_g2436(.A (inc_ADD_UNS_OP5492_3_n_2462), .B
       (csr_minstret[27]), .Q (n_7538));
  HAX1 inc_ADD_UNS_OP5492_3_g2437(.A (inc_ADD_UNS_OP5492_3_n_2468), .B
       (csr_minstret[35]), .S (n_7522), .CO
       (inc_ADD_UNS_OP5492_3_n_2459));
  HAX1 inc_ADD_UNS_OP5492_3_g2438(.A (inc_ADD_UNS_OP5492_3_n_2465), .B
       (csr_minstret[26]), .S (n_7540), .CO
       (inc_ADD_UNS_OP5492_3_n_2462));
  HAX1 inc_ADD_UNS_OP5492_3_g2439(.A (inc_ADD_UNS_OP5492_3_n_2474), .B
       (csr_minstret[25]), .S (n_7542), .CO
       (inc_ADD_UNS_OP5492_3_n_2465));
  EO2X1 inc_ADD_UNS_OP5492_3_g2440(.A (inc_ADD_UNS_OP5492_3_n_2472), .B
       (csr_minstret[34]), .Q (n_7524));
  AND5X1 inc_ADD_UNS_OP5492_3_g2441(.A (inc_ADD_UNS_OP5492_3_n_2490),
       .B (csr_minstret[31]), .C (csr_minstret[32]), .D
       (csr_minstret[33]), .E (csr_minstret[34]), .Q
       (inc_ADD_UNS_OP5492_3_n_2468));
  HAX1 inc_ADD_UNS_OP5492_3_g2442(.A (inc_ADD_UNS_OP5492_3_n_2476), .B
       (csr_minstret[33]), .S (n_7526), .CO
       (inc_ADD_UNS_OP5492_3_n_2472));
  HAX1 inc_ADD_UNS_OP5492_3_g2443(.A (inc_ADD_UNS_OP5492_3_n_2479), .B
       (csr_minstret[24]), .S (n_7544), .CO
       (inc_ADD_UNS_OP5492_3_n_2474));
  HAX1 inc_ADD_UNS_OP5492_3_g2444(.A (inc_ADD_UNS_OP5492_3_n_2480), .B
       (csr_minstret[32]), .S (n_7528), .CO
       (inc_ADD_UNS_OP5492_3_n_2476));
  HAX1 inc_ADD_UNS_OP5492_3_g2445(.A (inc_ADD_UNS_OP5492_3_n_2485), .B
       (csr_minstret[23]), .S (n_7546), .CO
       (inc_ADD_UNS_OP5492_3_n_2479));
  HAX2 inc_ADD_UNS_OP5492_3_g2446(.A (inc_ADD_UNS_OP5492_3_n_2490), .B
       (csr_minstret[31]), .S (n_7530), .CO
       (inc_ADD_UNS_OP5492_3_n_2480));
  HAX1 inc_ADD_UNS_OP5492_3_g2447(.A (inc_ADD_UNS_OP5492_3_n_2488), .B
       (csr_minstret[22]), .S (n_7548), .CO
       (inc_ADD_UNS_OP5492_3_n_2485));
  HAX1 inc_ADD_UNS_OP5492_3_g2448(.A (inc_ADD_UNS_OP5492_3_n_2497), .B
       (csr_minstret[21]), .S (n_7550), .CO
       (inc_ADD_UNS_OP5492_3_n_2488));
  EO2X1 inc_ADD_UNS_OP5492_3_g2449(.A (inc_ADD_UNS_OP5492_3_n_2493), .B
       (csr_minstret[30]), .Q (n_7532));
  AND3X4 inc_ADD_UNS_OP5492_3_g2450(.A (inc_ADD_UNS_OP5492_3_n_2498),
       .B (csr_minstret[29]), .C (csr_minstret[30]), .Q
       (inc_ADD_UNS_OP5492_3_n_2490));
  HAX1 inc_ADD_UNS_OP5492_3_g2451(.A (inc_ADD_UNS_OP5492_3_n_2498), .B
       (csr_minstret[29]), .S (n_7534), .CO
       (inc_ADD_UNS_OP5492_3_n_2493));
  HAX1 inc_ADD_UNS_OP5492_3_g2452(.A (inc_ADD_UNS_OP5492_3_n_2501), .B
       (csr_minstret[20]), .S (n_7552), .CO
       (inc_ADD_UNS_OP5492_3_n_2497));
  HAX2 inc_ADD_UNS_OP5492_3_g2453(.A (n_8600), .B (csr_minstret[28]),
       .S (n_7536), .CO (inc_ADD_UNS_OP5492_3_n_2498));
  HAX1 inc_ADD_UNS_OP5492_3_g2454(.A (inc_ADD_UNS_OP5492_3_n_2504), .B
       (csr_minstret[19]), .S (n_7554), .CO
       (inc_ADD_UNS_OP5492_3_n_2501));
  HAX2 inc_ADD_UNS_OP5492_3_g2456(.A (inc_ADD_UNS_OP5492_3_n_2507), .B
       (csr_minstret[18]), .S (n_7556), .CO
       (inc_ADD_UNS_OP5492_3_n_2504));
  HAX2 inc_ADD_UNS_OP5492_3_g2457(.A (inc_ADD_UNS_OP5492_3_n_2509), .B
       (csr_minstret[17]), .S (n_7558), .CO
       (inc_ADD_UNS_OP5492_3_n_2507));
  EO2X1 inc_ADD_UNS_OP5492_3_g2458(.A (inc_ADD_UNS_OP5492_3_n_2512), .B
       (csr_minstret[16]), .Q (n_7560));
  AND4X1 inc_ADD_UNS_OP5492_3_g2459(.A (inc_ADD_UNS_OP5492_3_n_2518),
       .B (csr_minstret[14]), .C (csr_minstret[15]), .D
       (csr_minstret[16]), .Q (inc_ADD_UNS_OP5492_3_n_2509));
  HAX1 inc_ADD_UNS_OP5492_3_g2460(.A (inc_ADD_UNS_OP5492_3_n_2515), .B
       (csr_minstret[15]), .S (n_7562), .CO
       (inc_ADD_UNS_OP5492_3_n_2512));
  HAX1 inc_ADD_UNS_OP5492_3_g2461(.A (inc_ADD_UNS_OP5492_3_n_2518), .B
       (csr_minstret[14]), .S (n_7564), .CO
       (inc_ADD_UNS_OP5492_3_n_2515));
  HAX1 inc_ADD_UNS_OP5492_3_g2462(.A (inc_ADD_UNS_OP5492_3_n_2521), .B
       (csr_minstret[13]), .S (n_7566), .CO
       (inc_ADD_UNS_OP5492_3_n_2518));
  HAX2 inc_ADD_UNS_OP5492_3_g2463(.A (inc_ADD_UNS_OP5492_3_n_2523), .B
       (csr_minstret[12]), .S (n_7568), .CO
       (inc_ADD_UNS_OP5492_3_n_2521));
  EO2X0 inc_ADD_UNS_OP5492_3_g2464(.A (inc_ADD_UNS_OP5492_3_n_2676), .B
       (csr_minstret[11]), .Q (n_7570));
  AND2X2 inc_ADD_UNS_OP5492_3_g2465(.A (inc_ADD_UNS_OP5492_3_n_2676),
       .B (csr_minstret[11]), .Q (inc_ADD_UNS_OP5492_3_n_2523));
  EO2X0 inc_ADD_UNS_OP5492_3_g2466(.A (inc_ADD_UNS_OP5492_3_n_2533), .B
       (csr_minstret[10]), .Q (n_7572));
  EO2X1 inc_ADD_UNS_OP5492_3_g2469(.A (inc_ADD_UNS_OP5492_3_n_2536), .B
       (csr_minstret[9]), .Q (n_7574));
  AND4X2 inc_ADD_UNS_OP5492_3_g2470(.A (inc_ADD_UNS_OP5492_3_n_2542),
       .B (csr_minstret[7]), .C (csr_minstret[8]), .D
       (csr_minstret[9]), .Q (inc_ADD_UNS_OP5492_3_n_2533));
  HAX1 inc_ADD_UNS_OP5492_3_g2471(.A (inc_ADD_UNS_OP5492_3_n_2539), .B
       (csr_minstret[8]), .S (n_7576), .CO
       (inc_ADD_UNS_OP5492_3_n_2536));
  HAX1 inc_ADD_UNS_OP5492_3_g2472(.A (inc_ADD_UNS_OP5492_3_n_2542), .B
       (csr_minstret[7]), .S (n_7578), .CO
       (inc_ADD_UNS_OP5492_3_n_2539));
  HAX2 inc_ADD_UNS_OP5492_3_g2473(.A (inc_ADD_UNS_OP5492_3_n_2545), .B
       (csr_minstret[6]), .S (n_7580), .CO
       (inc_ADD_UNS_OP5492_3_n_2542));
  EO2X0 inc_ADD_UNS_OP5492_3_g2474(.A (inc_ADD_UNS_OP5492_3_n_2553), .B
       (csr_minstret[5]), .Q (n_7582));
  AND2X4 inc_ADD_UNS_OP5492_3_g2475(.A (inc_ADD_UNS_OP5492_3_n_2553),
       .B (csr_minstret[5]), .Q (inc_ADD_UNS_OP5492_3_n_2545));
  EO2X1 inc_ADD_UNS_OP5492_3_g2476(.A (inc_ADD_UNS_OP5492_3_n_2551), .B
       (csr_minstret[3]), .Q (n_7586));
  HAX1 inc_ADD_UNS_OP5492_3_g2477(.A (inc_ADD_UNS_OP5492_3_n_2567), .B
       (csr_minstret[2]), .S (n_7588), .CO
       (inc_ADD_UNS_OP5492_3_n_2551));
  EN2X0 inc_ADD_UNS_OP5492_3_g2478(.A (inc_ADD_UNS_OP5492_3_n_2556), .B
       (csr_minstret[4]), .Q (n_7584));
  NO2I1X2 inc_ADD_UNS_OP5492_3_g2479(.B (inc_ADD_UNS_OP5492_3_n_2556),
       .AN (csr_minstret[4]), .Q (inc_ADD_UNS_OP5492_3_n_2553));
  NA3X2 inc_ADD_UNS_OP5492_3_g2480(.A (inc_ADD_UNS_OP5492_3_n_2567), .B
       (csr_minstret[2]), .C (csr_minstret[3]), .Q
       (inc_ADD_UNS_OP5492_3_n_2556));
  NO2I1X2 inc_ADD_UNS_OP5492_3_g2483(.B (inc_ADD_UNS_OP5492_3_n_2585),
       .AN (csr_minstret[1]), .Q (inc_ADD_UNS_OP5492_3_n_2567));
  AND5X1 inc_ADD_UNS_OP5492_3_g2485(.A (inc_ADD_UNS_OP5492_3_n_2580),
       .B (csr_minstret[45]), .C (csr_minstret[46]), .D
       (csr_minstret[50]), .E (csr_minstret[49]), .Q
       (inc_ADD_UNS_OP5492_3_n_2571));
  AND5X1 inc_ADD_UNS_OP5492_3_g2486(.A (csr_minstret[26]), .B
       (csr_minstret[27]), .C (csr_minstret[20]), .D
       (csr_minstret[19]), .E (csr_minstret[21]), .Q
       (inc_ADD_UNS_OP5492_3_n_2574));
  AND4X1 inc_ADD_UNS_OP5492_3_g2487(.A (csr_minstret[51]), .B
       (csr_minstret[47]), .C (csr_minstret[52]), .D
       (csr_minstret[48]), .Q (inc_ADD_UNS_OP5492_3_n_2580));
  EO2X1 inc_ADD_UNS_OP5492_3_g2488(.A (csr_minstret[0]), .B (n_7883),
       .Q (n_7592));
  NA2X2 inc_ADD_UNS_OP5492_3_g2489(.A (csr_minstret[0]), .B (n_7883),
       .Q (inc_ADD_UNS_OP5492_3_n_2585));
  INX1 inc_ADD_UNS_OP5492_3_g2495(.A (csr_minstret[55]), .Q
       (inc_ADD_UNS_OP5492_3_n_2608));
  INX1 inc_ADD_UNS_OP5492_3_g2497(.A (csr_minstret[45]), .Q
       (inc_ADD_UNS_OP5492_3_n_2613));
  INX1 inc_ADD_UNS_OP5492_3_g2498(.A (csr_minstret[50]), .Q
       (inc_ADD_UNS_OP5492_3_n_2615));
  INX1 inc_ADD_UNS_OP5492_3_g2504(.A (csr_minstret[61]), .Q
       (inc_ADD_UNS_OP5492_3_n_2647));
  INX1 inc_ADD_UNS_OP5492_3_g2505(.A (csr_minstret[59]), .Q
       (inc_ADD_UNS_OP5492_3_n_2649));
  INX1 inc_ADD_UNS_OP5492_3_g2507(.A (csr_minstret[57]), .Q
       (inc_ADD_UNS_OP5492_3_n_2656));
  EO2X1 inc_ADD_UNS_OP5492_3_g2(.A (inc_ADD_UNS_OP5492_3_n_2339), .B
       (csr_minstret[62]), .Q (n_7468));
  EO2X1 inc_ADD_UNS_OP5492_3_g2510(.A (inc_ADD_UNS_OP5492_3_n_2350), .B
       (csr_minstret[60]), .Q (n_7472));
  EO2X1 inc_ADD_UNS_OP5492_3_g2511(.A (inc_ADD_UNS_OP5492_3_n_2366), .B
       (csr_minstret[51]), .Q (n_7490));
  EO2X1 inc_ADD_UNS_OP5492_3_g2512(.A (inc_ADD_UNS_OP5492_3_n_2371), .B
       (csr_minstret[58]), .Q (n_7476));
  EO2X1 inc_ADD_UNS_OP5492_3_g2513(.A (inc_ADD_UNS_OP5492_3_n_2380), .B
       (csr_minstret[49]), .Q (n_7494));
  EO2X1 inc_ADD_UNS_OP5492_3_g2514(.A (inc_ADD_UNS_OP5492_3_n_2388), .B
       (csr_minstret[56]), .Q (n_7480));
  EO2X1 inc_ADD_UNS_OP5492_3_g2515(.A (inc_ADD_UNS_OP5492_3_n_2409), .B
       (csr_minstret[54]), .Q (n_7484));
  EO2X1 inc_ADD_UNS_OP5492_3_g2516(.A (inc_ADD_UNS_OP5492_3_n_2413), .B
       (csr_minstret[46]), .Q (n_7500));
  NA2I1X1 inc_ADD_UNS_OP5492_3_g2517(.B (inc_ADD_UNS_OP5492_3_n_2571),
       .AN (inc_ADD_UNS_OP5492_3_n_2419), .Q
       (inc_ADD_UNS_OP5492_3_n_2675));
  AND2X1 inc_ADD_UNS_OP5492_3_g2518(.A (inc_ADD_UNS_OP5492_3_n_2533),
       .B (csr_minstret[10]), .Q (inc_ADD_UNS_OP5492_3_n_2676));
  EN2X0 inc_ADD_UNS_OP5492_3_g2519(.A (inc_ADD_UNS_OP5492_3_n_2585), .B
       (csr_minstret[1]), .Q (n_7590));
  EO2X1 inc_ADD_UNS_OP5492_3_g2520(.A (inc_ADD_UNS_OP5492_3_n_2439), .B
       (csr_minstret[41]), .Q (n_7510));
  EN2X1 inc_ADD_UNS_OP5492_3_g2521(.A (inc_ADD_UNS_OP5492_3_n_2356), .B
       (csr_minstret[52]), .Q (n_7488));
  EN2X1 inc_ADD_UNS_OP5492_3_g2522(.A (inc_ADD_UNS_OP5492_3_n_2430), .B
       (csr_minstret[43]), .Q (n_7506));
  EN2X1 inc_ADD_UNS_OP5492_3_g2523(.A (inc_ADD_UNS_OP5492_3_n_2427), .B
       (csr_minstret[44]), .Q (n_7504));
  EN2X1 inc_ADD_UNS_OP5492_3_g2524(.A (inc_ADD_UNS_OP5492_3_n_2675), .B
       (csr_minstret[53]), .Q (n_7486));
  EO2X1 add_1545_30_g1380(.A (add_1545_30_n_811), .B (csr_mtvec[19]),
       .Q (n_7841));
  EO2X1 add_1545_30_g1381(.A (add_1545_30_n_814), .B (csr_mtvec[15]),
       .Q (n_7845));
  HAX1 add_1545_30_g1382(.A (add_1545_30_n_821), .B (csr_mtvec[18]), .S
       (n_7842), .CO (add_1545_30_n_811));
  EO2X1 add_1545_30_g1383(.A (add_1545_30_n_816), .B (csr_mtvec[11]),
       .Q (n_7849));
  HAX1 add_1545_30_g1384(.A (add_1545_30_n_827), .B (csr_mtvec[14]), .S
       (n_7846), .CO (add_1545_30_n_814));
  HAX1 add_1545_30_g1385(.A (add_1545_30_n_835), .B (csr_mtvec[10]), .S
       (n_7850), .CO (add_1545_30_n_816));
  EO2X1 add_1545_30_g1386(.A (add_1545_30_n_825), .B (csr_mtvec[27]),
       .Q (n_7833));
  EO2X1 add_1545_30_g1387(.A (add_1545_30_n_831), .B (csr_mtvec[31]),
       .Q (n_7829));
  EO2X1 add_1545_30_g1388(.A (add_1545_30_n_829), .B (csr_mtvec[23]),
       .Q (n_7837));
  HAX1 add_1545_30_g1389(.A (add_1545_30_n_840), .B (csr_mtvec[17]), .S
       (n_7843), .CO (add_1545_30_n_821));
  EO2X1 add_1545_30_g1390(.A (add_1545_30_n_833), .B (csr_mtvec[25]),
       .Q (n_7835));
  EO2X1 add_1545_30_g1391(.A (add_1545_30_n_837), .B (csr_mtvec[21]),
       .Q (n_7839));
  HAX1 add_1545_30_g1392(.A (add_1545_30_n_847), .B (csr_mtvec[26]), .S
       (n_7834), .CO (add_1545_30_n_825));
  HAX1 add_1545_30_g1393(.A (add_1545_30_n_843), .B (csr_mtvec[13]), .S
       (n_7847), .CO (add_1545_30_n_827));
  HAX1 add_1545_30_g1394(.A (add_1545_30_n_851), .B (csr_mtvec[22]), .S
       (n_7838), .CO (add_1545_30_n_829));
  HAX1 add_1545_30_g1395(.A (add_1545_30_n_848), .B (csr_mtvec[30]), .S
       (n_7830), .CO (add_1545_30_n_831));
  HAX1 add_1545_30_g1396(.A (add_1545_30_n_858), .B (csr_mtvec[24]), .S
       (n_7836), .CO (add_1545_30_n_833));
  HAX1 add_1545_30_g1397(.A (add_1545_30_n_854), .B (csr_mtvec[9]), .S
       (n_7851), .CO (add_1545_30_n_835));
  HAX1 add_1545_30_g1398(.A (add_1545_30_n_860), .B (csr_mtvec[20]), .S
       (n_7840), .CO (add_1545_30_n_837));
  EN2X1 add_1545_30_g1399(.A (add_1545_30_n_844), .B (csr_mtvec[29]),
       .Q (n_7831));
  HAX1 add_1545_30_g1400(.A (add_1545_30_n_861), .B (csr_mtvec[16]), .S
       (n_7844), .CO (add_1545_30_n_840));
  EN2X0 add_1545_30_g1401(.A (add_1545_30_n_855), .B (csr_mtvec[28]),
       .Q (n_7832));
  HAX1 add_1545_30_g1402(.A (add_1545_30_n_867), .B (csr_mtvec[12]), .S
       (n_7848), .CO (add_1545_30_n_843));
  NA3X1 add_1545_30_g1403(.A (add_1545_30_n_858), .B
       (add_1545_30_n_888), .C (csr_mtvec[28]), .Q (add_1545_30_n_844));
  NO2I1X1 add_1545_30_g1404(.B (add_1545_30_n_904), .AN
       (add_1545_30_n_858), .Q (add_1545_30_n_847));
  NO3I2X1 add_1545_30_g1405(.C (add_1545_30_n_855), .AN
       (csr_mtvec[29]), .BN (csr_mtvec[28]), .Q (add_1545_30_n_848));
  NO2I1X1 add_1545_30_g1406(.B (add_1545_30_n_898), .AN
       (add_1545_30_n_860), .Q (add_1545_30_n_851));
  HAX1 add_1545_30_g1407(.A (add_1545_30_n_873), .B (csr_mtvec[8]), .S
       (n_7852), .CO (add_1545_30_n_854));
  NA3X1 add_1545_30_g1408(.A (add_1545_30_n_861), .B
       (add_1545_30_n_883), .C (add_1545_30_n_888), .Q
       (add_1545_30_n_855));
  AND2X1 add_1545_30_g1409(.A (add_1545_30_n_861), .B
       (add_1545_30_n_883), .Q (add_1545_30_n_858));
  AND2X1 add_1545_30_g1410(.A (add_1545_30_n_861), .B
       (add_1545_30_n_892), .Q (add_1545_30_n_860));
  AND5X1 add_1545_30_g1411(.A (add_1545_30_n_867), .B (csr_mtvec[12]),
       .C (csr_mtvec[13]), .D (csr_mtvec[15]), .E (csr_mtvec[14]), .Q
       (add_1545_30_n_861));
  AND5X1 add_1545_30_g1412(.A (add_1545_30_n_873), .B (csr_mtvec[8]),
       .C (csr_mtvec[9]), .D (csr_mtvec[11]), .E (csr_mtvec[10]), .Q
       (add_1545_30_n_867));
  HAX1 add_1545_30_g1413(.A (add_1545_30_n_876), .B (csr_mtvec[7]), .S
       (n_7853), .CO (add_1545_30_n_873));
  FAX1 add_1545_30_g1414(.A (csr_mtvec[6]), .B (csr_mcause_code[4]),
       .CI (add_1545_30_n_878), .S (n_7854), .CO (add_1545_30_n_876));
  FAX1 add_1545_30_g1415(.A (csr_mtvec[5]), .B (csr_mcause_code[3]),
       .CI (add_1545_30_n_880), .S (n_7855), .CO (add_1545_30_n_878));
  FAX1 add_1545_30_g1416(.A (csr_mtvec[4]), .B (csr_mcause_code[2]),
       .CI (add_1545_30_n_882), .S (n_7856), .CO (add_1545_30_n_880));
  FAX1 add_1545_30_g1417(.A (csr_mtvec[3]), .B (csr_mcause_code[1]),
       .CI (n_8665), .S (n_7857), .CO (add_1545_30_n_882));
  NO3I1X1 add_1545_30_g1418(.B (add_1545_30_n_898), .C
       (add_1545_30_n_901), .AN (add_1545_30_n_892), .Q
       (add_1545_30_n_883));
  NO3I2X1 add_1545_30_g1420(.C (add_1545_30_n_904), .AN
       (csr_mtvec[27]), .BN (csr_mtvec[26]), .Q (add_1545_30_n_888));
  AND4X1 add_1545_30_g1421(.A (csr_mtvec[18]), .B (csr_mtvec[16]), .C
       (csr_mtvec[19]), .D (csr_mtvec[17]), .Q (add_1545_30_n_892));
  NA2X1 add_1545_30_g1423(.A (csr_mtvec[20]), .B (csr_mtvec[21]), .Q
       (add_1545_30_n_898));
  NA2X1 add_1545_30_g1424(.A (csr_mtvec[22]), .B (csr_mtvec[23]), .Q
       (add_1545_30_n_901));
  NA2X1 add_1545_30_g1425(.A (csr_mtvec[24]), .B (csr_mtvec[25]), .Q
       (add_1545_30_n_904));
  EO2X1 add_459_21_g964(.A (add_459_21_n_642), .B
       (program_counter[27]), .Q (n_7952));
  EO2X1 add_459_21_g965(.A (add_459_21_n_645), .B
       (program_counter[23]), .Q (n_7947));
  HAX1 add_459_21_g966(.A (add_459_21_n_652), .B (program_counter[26]),
       .S (n_7951), .CO (add_459_21_n_642));
  EO2X1 add_459_21_g967(.A (add_459_21_n_648), .B
       (program_counter[19]), .Q (n_7943));
  HAX1 add_459_21_g968(.A (add_459_21_n_660), .B (program_counter[22]),
       .S (n_7946), .CO (add_459_21_n_645));
  EO2X1 add_459_21_g969(.A (add_459_21_n_654), .B
       (program_counter[15]), .Q (n_7939));
  HAX1 add_459_21_g970(.A (add_459_21_n_664), .B (program_counter[18]),
       .S (n_7942), .CO (add_459_21_n_648));
  EO2X1 add_459_21_g971(.A (add_459_21_n_658), .B
       (program_counter[31]), .Q (n_7956));
  EO2X1 add_459_21_g972(.A (add_459_21_n_662), .B
       (program_counter[11]), .Q (n_7935));
  HAX1 add_459_21_g973(.A (add_459_21_n_670), .B (program_counter[25]),
       .S (n_7950), .CO (add_459_21_n_652));
  HAX1 add_459_21_g974(.A (add_459_21_n_672), .B (program_counter[14]),
       .S (n_7938), .CO (add_459_21_n_654));
  EO2X1 add_459_21_g975(.A (add_459_21_n_668), .B
       (program_counter[29]), .Q (n_7954));
  EO2X1 add_459_21_g976(.A (add_459_21_n_666), .B (program_counter[7]),
       .Q (n_7931));
  HAX1 add_459_21_g977(.A (add_459_21_n_677), .B (program_counter[30]),
       .S (n_7955), .CO (add_459_21_n_658));
  HAX1 add_459_21_g978(.A (add_459_21_n_676), .B (program_counter[21]),
       .S (n_7945), .CO (add_459_21_n_660));
  HAX1 add_459_21_g979(.A (add_459_21_n_674), .B (program_counter[10]),
       .S (n_7934), .CO (add_459_21_n_662));
  HAX1 add_459_21_g980(.A (add_459_21_n_684), .B (program_counter[17]),
       .S (n_7941), .CO (add_459_21_n_664));
  HAX1 add_459_21_g981(.A (add_459_21_n_682), .B (program_counter[6]),
       .S (n_7930), .CO (add_459_21_n_666));
  HAX1 add_459_21_g982(.A (add_459_21_n_685), .B (program_counter[28]),
       .S (n_7953), .CO (add_459_21_n_668));
  HAX1 add_459_21_g983(.A (add_459_21_n_693), .B (program_counter[24]),
       .S (n_7948), .CO (add_459_21_n_670));
  HAX1 add_459_21_g984(.A (add_459_21_n_692), .B (program_counter[13]),
       .S (n_7937), .CO (add_459_21_n_672));
  HAX1 add_459_21_g985(.A (add_459_21_n_700), .B (program_counter[9]),
       .S (n_7933), .CO (add_459_21_n_674));
  HAX1 add_459_21_g986(.A (add_459_21_n_701), .B (program_counter[20]),
       .S (n_7944), .CO (add_459_21_n_676));
  AND3X1 add_459_21_g987(.A (add_459_21_n_685), .B
       (program_counter[28]), .C (program_counter[29]), .Q
       (add_459_21_n_677));
  HAX1 add_459_21_g988(.A (add_459_21_n_708), .B (program_counter[5]),
       .S (n_7929), .CO (add_459_21_n_682));
  HAX1 add_459_21_g989(.A (add_459_21_n_709), .B (program_counter[16]),
       .S (n_7940), .CO (add_459_21_n_684));
  AND5X1 add_459_21_g990(.A (add_459_21_n_693), .B
       (program_counter[24]), .C (program_counter[25]), .D
       (program_counter[27]), .E (program_counter[26]), .Q
       (add_459_21_n_685));
  HAX1 add_459_21_g991(.A (add_459_21_n_715), .B (program_counter[12]),
       .S (n_7936), .CO (add_459_21_n_692));
  AND5X1 add_459_21_g992(.A (add_459_21_n_701), .B
       (program_counter[20]), .C (program_counter[21]), .D
       (program_counter[23]), .E (program_counter[22]), .Q
       (add_459_21_n_693));
  HAX1 add_459_21_g993(.A (add_459_21_n_721), .B (program_counter[8]),
       .S (n_7932), .CO (add_459_21_n_700));
  AND5X1 add_459_21_g994(.A (add_459_21_n_709), .B
       (program_counter[16]), .C (program_counter[17]), .D
       (program_counter[19]), .E (program_counter[18]), .Q
       (add_459_21_n_701));
  HAX1 add_459_21_g995(.A (add_459_21_n_727), .B (program_counter[4]),
       .S (n_7927), .CO (add_459_21_n_708));
  AND5X1 add_459_21_g996(.A (add_459_21_n_715), .B
       (program_counter[12]), .C (program_counter[13]), .D
       (program_counter[15]), .E (program_counter[14]), .Q
       (add_459_21_n_709));
  AND5X1 add_459_21_g997(.A (add_459_21_n_721), .B
       (program_counter[8]), .C (program_counter[9]), .D
       (program_counter[11]), .E (program_counter[10]), .Q
       (add_459_21_n_715));
  AND5X1 add_459_21_g998(.A (add_459_21_n_727), .B
       (program_counter[4]), .C (program_counter[5]), .D
       (program_counter[7]), .E (program_counter[6]), .Q
       (add_459_21_n_721));
  HAX1 add_459_21_g999(.A (program_counter[2]), .B
       (program_counter[3]), .S (n_7926), .CO (add_459_21_n_727));
  INX2 g92631(.A (n_4673), .Q (n_4677));
  MU2X1 g92638(.S (alu_2nd_operand[13]), .IN0
       (alu_operation_code_39112), .IN1 (n_2326), .Q (n_8311));
  EN2X1 g92639(.A (n_4224), .B (alu_operation_code_39112), .Q (n_8312));
  EN2X1 g92640(.A (n_4225), .B (alu_operation_code_39112), .Q (n_8313));
  EN2X1 g92641(.A (n_8497), .B (alu_operation_code_39112), .Q (n_8314));
  MU2X1 g92642(.S (n_8495), .IN0 (alu_operation_code_39112), .IN1
       (n_2326), .Q (n_8315));
  EN2X1 g92643(.A (n_2326), .B (n_8677), .Q (n_8316));
  MU2X1 g92644(.S (n_2258), .IN0 (n_7671), .IN1 (n_4151), .Q (n_8317));
  MU2X1 g3(.S (add_463_14_n_836), .IN0 (add_463_14_n_748), .IN1
       (add_463_14_n_749), .Q (n_8318));
  NA2X2 g92646(.A (n_8320), .B (n_175), .Q (n_8321));
  EN2X1 g92647(.A (inc_add_1343_59_4_n_3386), .B
       (inc_add_1343_59_4_n_3769), .Q (n_8320));
  NA2X2 g92648(.A (n_8322), .B (n_175), .Q (n_8323));
  EN2X1 g92649(.A (inc_add_1343_59_4_n_3413), .B
       (inc_add_1343_59_4_n_3749), .Q (n_8322));
  NA2X2 g92652(.A (n_8326), .B (n_159), .Q (n_8327));
  EN2X1 g92653(.A (inc_ADD_UNS_OP_5_n_3370), .B
       (inc_ADD_UNS_OP_5_n_3735), .Q (n_8326));
  NA2X2 g92654(.A (n_8364), .B (n_159), .Q (n_8329));
  NA2X1 g92656(.A (n_8330), .B (n_159), .Q (n_8331));
  EO2X1 g92657(.A (n_8596), .B (csr_minstret[35]), .Q (n_8330));
  NA2X1 g92658(.A (n_8332), .B (n_159), .Q (n_8333));
  EN2X1 g92659(.A (inc_ADD_UNS_OP_5_n_3400), .B
       (inc_ADD_UNS_OP_5_n_3793), .Q (n_8332));
  NA2X1 g92660(.A (n_8363), .B (n_159), .Q (n_8335));
  NA2X1 g92662(.A (n_8362), .B (n_159), .Q (n_8337));
  NA2X1 g92664(.A (n_8338), .B (n_159), .Q (n_8339));
  EN2X1 g92665(.A (inc_ADD_UNS_OP_5_n_3392), .B
       (inc_ADD_UNS_OP_5_n_3782), .Q (n_8338));
  AN21X1 g92666(.A (n_7370), .B (n_1082), .C (n_1081), .Q (n_8340));
  AN21X1 g92667(.A (add_463_14_n_800), .B (n_8341), .C
       (add_463_14_n_776), .Q (n_8342));
  AO21X1 g92668(.A (add_463_14_n_760), .B (add_463_14_n_646), .C
       (add_463_14_n_699), .Q (n_8341));
  AN21X1 g92669(.A (add_464_21_n_811), .B (n_8343), .C
       (add_464_21_n_752), .Q (n_8344));
  AO21X1 g92670(.A (add_464_21_n_708), .B (add_464_21_n_637), .C
       (add_464_21_n_686), .Q (n_8343));
  AN21X1 g92671(.A (add_464_21_n_812), .B (n_8345), .C
       (add_464_21_n_750), .Q (n_8346));
  AO21X1 g92672(.A (add_464_21_n_730), .B (add_464_21_n_637), .C
       (add_464_21_n_701), .Q (n_8345));
  AN21X1 g92673(.A (add_464_21_n_878), .B (n_8347), .C
       (add_464_21_n_863), .Q (n_8348));
  AO21X1 g92674(.A (add_464_21_n_768), .B (add_464_21_n_637), .C
       (add_464_21_n_729), .Q (n_8347));
  EO2X1 g92675(.A (inc_ADD_UNS_OP_5_n_3411), .B (n_7377), .Q (n_8349));
  EN2X1 g92676(.A (inc_ADD_UNS_OP5491_6_n_2366), .B
       (inc_add_1345_58_1_n_3455), .Q (n_8350));
  EN2X1 g92677(.A (inc_add_1347_34_2_n_2311), .B (csr_mcycle[63]), .Q
       (n_8351));
  EN2X1 g92678(.A (inc_add_1347_34_2_n_2316), .B (csr_mcycle[55]), .Q
       (n_8352));
  EN2X1 g92679(.A (inc_ADD_UNS_OP5492_3_n_2334), .B (csr_minstret[63]),
       .Q (n_8353));
  OR2X4 g92680(.A (n_2345), .B (n_2672), .Q (n_8354));
  AND2X4 g92681(.A (n_906), .B (n_905), .Q (n_8355));
  NA3I2X2 g92684(.C (n_2495), .AN (n_2625), .BN (n_2263), .Q (n_8358));
  OR2X4 g92685(.A (n_8481), .B (instruction[28]), .Q (n_8359));
  NA2I1X2 g92686(.B (n_2477), .AN (n_2306), .Q (n_8360));
  NO2I1X4 g92687(.B (n_8588), .AN (n_178), .Q (n_8361));
  EO2X1 g92688(.A (inc_ADD_UNS_OP_5_n_3415), .B
       (inc_ADD_UNS_OP_5_n_3792), .Q (n_8362));
  EO2X1 g92689(.A (inc_ADD_UNS_OP_5_n_3445), .B
       (inc_ADD_UNS_OP_5_n_3785), .Q (n_8363));
  EO2X1 g92690(.A (inc_ADD_UNS_OP_5_n_3421), .B (csr_minstret[33]), .Q
       (n_8364));
  NA3I2X1 g92691(.C (n_2243), .AN (n_4369), .BN (n_8218), .Q (n_8365));
  NA5I1X4 g92692(.B (n_6060), .C (n_5995), .D (n_5371), .E (n_5357),
       .AN (n_8453), .Q (n_8366));
  NO3I2X2 g92696(.C (n_8663), .AN (n_5808), .BN (n_8617), .Q (n_8370));
  NA3I2X1 g92697(.C (n_8418), .AN (n_5728), .BN (n_5711), .Q (n_8371));
  NA3X2 g92698(.A (n_5721), .B (n_5665), .C (n_8416), .Q (n_8372));
  NA3I2X1 g92701(.C (n_8432), .AN (n_5581), .BN (n_5652), .Q (n_8375));
  NA3I2X1 g92702(.C (n_8425), .AN (n_5623), .BN (n_5693), .Q (n_8376));
  NA3I2X2 g92703(.C (n_4522), .AN (n_4998), .BN (n_5684), .Q (n_8377));
  NA3X1 g92704(.A (n_8420), .B (n_5561), .C (n_5567), .Q (n_8378));
  NA3I2X2 g92705(.C (n_8433), .AN (n_5578), .BN (n_5651), .Q (n_8379));
  NA3X1 g92708(.A (n_5878), .B (n_5550), .C (n_5556), .Q (n_8382));
  NA3I2X2 g92709(.C (n_8696), .AN (n_5555), .BN (n_5549), .Q (n_8383));
  NA3X2 g92712(.A (n_5535), .B (n_8457), .C (n_8488), .Q (n_8386));
  NA3I2X2 g92713(.C (n_8616), .AN (n_5495), .BN (n_5511), .Q (n_8387));
  NA3I2X1 g92714(.C (n_8697), .AN (n_5494), .BN (n_5509), .Q (n_8388));
  NA3X1 g92717(.A (n_5823), .B (n_5432), .C (n_5445), .Q (n_8391));
  NA3I2X2 g92718(.C (n_4517), .AN (n_5458), .BN (n_5443), .Q (n_8392));
  NA3I2X2 g92720(.C (n_5807), .AN (n_5451), .BN (n_5435), .Q (n_8394));
  NA3I2X2 g92722(.C (n_5805), .AN (n_5430), .BN (n_8467), .Q (n_8396));
  NO3I1X1 g92723(.B (n_5410), .C (n_8469), .AN (n_8451), .Q (n_8397));
  NO5X4 g92726(.A (n_5768), .B (n_4932), .C (n_4933), .D (n_4964), .E
       (n_4965), .Q (n_8400));
  NO6X4 g92727(.A (n_4920), .B (n_4913), .C (n_4952), .D (n_4938), .E
       (n_8470), .F (n_5383), .Q (n_8401));
  NO5X4 g92728(.A (n_5761), .B (n_4912), .C (n_4910), .D (n_4945), .E
       (n_4939), .Q (n_8402));
  NO5X4 g92729(.A (n_5774), .B (n_4969), .C (n_4966), .D (n_4982), .E
       (n_4983), .Q (n_8403));
  NO6X4 g92731(.A (n_4854), .B (n_4855), .C (n_4856), .D (n_4857), .E
       (n_8472), .F (n_8471), .Q (n_8405));
  AN221X1 g92737(.A (n_4901), .B (n_6371), .C (n_4899), .D (n_6367), .E
       (n_5713), .Q (n_8411));
  AN221X1 g92738(.A (n_4893), .B (n_6945), .C (n_4891), .D (n_6941), .E
       (n_5707), .Q (n_8412));
  AN222X1 g92739(.A (n_4741), .B (n_7218), .C (n_4903), .D (n_7223), .E
       (n_4861), .F (n_7219), .Q (n_8413));
  AN222X1 g92740(.A (n_4741), .B (n_6412), .C (n_4903), .D (n_6417), .E
       (n_4861), .F (n_6413), .Q (n_8414));
  AN222X1 g92741(.A (n_4741), .B (n_6939), .C (n_4903), .D (n_6944), .E
       (n_4861), .F (n_6940), .Q (n_8415));
  AN221X1 g92742(.A (n_4897), .B (n_6988), .C (n_4895), .D (n_6992), .E
       (n_5729), .Q (n_8416));
  AN221X1 g92743(.A (n_4893), .B (n_6976), .C (n_4891), .D (n_6972), .E
       (n_5678), .Q (n_8417));
  AN221X1 g92744(.A (n_4508), .B (n_6906), .C (n_4503), .D (n_6907), .E
       (n_5720), .Q (n_8418));
  AN221X1 g92745(.A (n_4903), .B (n_6355), .C (n_4861), .D (n_6351), .E
       (n_4997), .Q (n_8419));
  AN222X1 g92746(.A (n_4741), .B (n_6877), .C (n_4903), .D (n_6882), .E
       (n_4861), .F (n_6878), .Q (n_8420));
  AN221X1 g92747(.A (n_4873), .B (n_6313), .C (n_4882), .D (n_6314), .E
       (n_5677), .Q (n_8421));
  AN221X1 g92748(.A (n_4873), .B (n_6561), .C (n_4882), .D (n_6562), .E
       (n_5674), .Q (n_8422));
  AN221X1 g92749(.A (n_4901), .B (n_7115), .C (n_4899), .D (n_7111), .E
       (n_5671), .Q (n_8423));
  AN221X1 g92750(.A (n_4866), .B (n_6950), .C (n_4497), .D (n_6951), .E
       (n_5612), .Q (n_8424));
  AN221X1 g92751(.A (n_4508), .B (n_6286), .C (n_4503), .D (n_6287), .E
       (n_5675), .Q (n_8425));
  AN221X1 g92752(.A (n_4508), .B (n_6875), .C (n_4502), .D (n_6876), .E
       (n_5649), .Q (n_8426));
  AN221X1 g92753(.A (n_4883), .B (n_6841), .C (n_4873), .D (n_6840), .E
       (n_5648), .Q (n_8427));
  AN221X1 g92754(.A (n_4876), .B (n_6845), .C (n_4508), .D (n_6844), .E
       (n_5656), .Q (n_8428));
  AN221X1 g92755(.A (n_4508), .B (n_7185), .C (n_4876), .D (n_7186), .E
       (n_5647), .Q (n_8429));
  AN221X1 g92756(.A (n_4901), .B (n_7146), .C (n_4899), .D (n_7142), .E
       (n_5646), .Q (n_8430));
  AN221X1 g92758(.A (n_4508), .B (n_7030), .C (n_4503), .D (n_7031), .E
       (n_5644), .Q (n_8432));
  AN221X1 g92759(.A (n_4897), .B (n_6337), .C (n_4895), .D (n_6341), .E
       (n_5579), .Q (n_8433));
  AN221X1 g92760(.A (n_4883), .B (n_6934), .C (n_4452), .D (n_6933), .E
       (n_5658), .Q (n_8434));
  AN221X1 g92761(.A (n_4878), .B (n_6890), .C (n_4506), .D (n_6891), .E
       (n_5576), .Q (n_8435));
  AN221X1 g92762(.A (n_4893), .B (n_6821), .C (n_4891), .D (n_6817), .E
       (n_5609), .Q (n_8436));
  AN221X1 g92764(.A (n_4893), .B (n_6294), .C (n_4891), .D (n_6290), .E
       (n_5546), .Q (n_8438));
  AN221X1 g92765(.A (n_4893), .B (n_6263), .C (n_4891), .D (n_6259), .E
       (n_5545), .Q (n_8439));
  AN221X1 g92766(.A (n_4866), .B (n_6981), .C (n_4498), .D (n_6982), .E
       (n_5562), .Q (n_8440));
  AN221X1 g92767(.A (n_4506), .B (n_6550), .C (n_4878), .D (n_6549), .E
       (n_5544), .Q (n_8441));
  AN221X1 g92768(.A (n_4893), .B (n_6325), .C (n_4891), .D (n_6321), .E
       (n_5523), .Q (n_8442));
  AN221X1 g92772(.A (n_4506), .B (n_6767), .C (n_4878), .D (n_6766), .E
       (n_5501), .Q (n_8446));
  NO3I1X2 g92776(.B (n_5043), .C (n_5044), .AN (n_5423), .Q (n_8450));
  AN211X1 g92777(.A (n_4481), .B (n_7233), .C (n_8468), .D (n_5034), .Q
       (n_8451));
  NA3I2X1 g92779(.C (n_5358), .AN (n_4831), .BN (n_4832), .Q (n_8453));
  NA3I2X1 g92780(.C (n_5342), .AN (n_4782), .BN (n_4787), .Q (n_8454));
  AO22X1 g92782(.A (n_4876), .B (n_6938), .C (n_4508), .D (n_6937), .Q
       (n_8456));
  AN21X1 g92783(.A (n_4508), .B (n_7061), .C (n_5190), .Q (n_8457));
  AN21X1 g92784(.A (n_4508), .B (n_6751), .C (n_5159), .Q (n_8458));
  AO22X2 g92785(.A (n_4893), .B (n_6573), .C (n_4891), .D (n_6569), .Q
       (n_8459));
  AO22X2 g92786(.A (n_4498), .B (n_6703), .C (n_4499), .D (n_6702), .Q
       (n_8460));
  AO22X2 g92787(.A (n_4868), .B (n_6570), .C (n_4870), .D (n_6571), .Q
       (n_8461));
  AO22X2 g92788(.A (n_4499), .B (n_6578), .C (n_4498), .D (n_6579), .Q
       (n_8462));
  AN21X1 g92789(.A (n_4893), .B (n_6635), .C (n_5123), .Q (n_8463));
  AO22X2 g92790(.A (n_4508), .B (n_6503), .C (n_4503), .D (n_6504), .Q
       (n_8464));
  AN22X1 g92791(.A (n_4878), .B (n_6642), .C (n_4506), .D (n_6643), .Q
       (n_8465));
  AO22X2 g92793(.A (n_4889), .B (n_6483), .C (n_4884), .D (n_6484), .Q
       (n_8467));
  AO22X1 g92794(.A (n_4489), .B (n_7241), .C (n_4738), .D (n_7242), .Q
       (n_8468));
  AO22X1 g92795(.A (n_4745), .B (n_7237), .C (n_4488), .D (n_7238), .Q
       (n_8469));
  AO22X1 g92796(.A (n_4481), .B (n_7171), .C (n_4491), .D (n_7172), .Q
       (n_8470));
  AO22X1 g92797(.A (n_4481), .B (n_6334), .C (n_4491), .D (n_6335), .Q
       (n_8471));
  AO22X1 g92798(.A (n_4489), .B (n_6342), .C (n_4738), .D (n_6343), .Q
       (n_8472));
  AN21X1 g92799(.A (n_4484), .B (n_6749), .C (n_4803), .Q (n_8473));
  AN21X1 g92800(.A (n_4745), .B (n_6710), .C (n_4795), .Q (n_8474));
  AN21X1 g92801(.A (n_4484), .B (n_6718), .C (n_4800), .Q (n_8475));
  AN21X1 g92802(.A (n_4484), .B (n_6687), .C (n_4860), .Q (n_8476));
  AN21X1 g92803(.A (n_4492), .B (n_6730), .C (n_4789), .Q (n_8477));
  AO22X1 g92804(.A (n_4745), .B (n_6493), .C (n_4488), .D (n_6494), .Q
       (n_8478));
  OA21X2 g92805(.A (n_4724), .B (jal_type), .C (n_4708), .Q (n_8479));
  AO22X2 g92806(.A (n_8224), .B (prev_instruction[27]), .C (n_4585), .D
       (read_data[27]), .Q (n_8480));
  AO22X2 g92807(.A (n_4465), .B (prev_instruction[29]), .C (n_4467), .D
       (read_data[29]), .Q (n_8481));
  AO22X4 g92808(.A (n_8224), .B (prev_instruction[31]), .C (n_4585), .D
       (read_data[31]), .Q (n_8482));
  AO22X4 g92810(.A (n_8224), .B (prev_instruction[30]), .C (n_4585), .D
       (read_data[30]), .Q (n_8484));
  AO22X2 g92811(.A (n_4585), .B (read_data[25]), .C (n_4465), .D
       (prev_instruction[25]), .Q (n_8485));
  AO22X2 g92812(.A (n_8224), .B (prev_instruction[26]), .C (n_4467), .D
       (read_data[26]), .Q (n_8486));
  AO22X4 g92813(.A (n_8224), .B (prev_instruction[13]), .C (n_4467), .D
       (read_data[13]), .Q (n_8487));
  NO3I1X2 g92814(.B (n_5199), .C (n_5200), .AN (n_5538), .Q (n_8488));
  OA22X2 g92815(.A (n_4264), .B (n_4247), .C (n_4246), .D (n_4181), .Q
       (n_8489));
  AO22X2 g92816(.A (alu_2nd_operand[14]), .B (n_2326), .C (n_4243), .D
       (alu_operation_code_39112), .Q (n_8490));
  AO22X2 g92817(.A (alu_2nd_operand[20]), .B (n_2326), .C (n_4223), .D
       (alu_operation_code_39112), .Q (n_8491));
  NO3X2 g92818(.A (n_4244), .B (n_4208), .C (n_2379), .Q (n_8492));
  AO22X2 g92819(.A (n_4153), .B (n_6141), .C (n_4141), .D
       (\rs1_data[19]_39596 ), .Q (n_8493));
  OA22X2 g92820(.A (n_4131), .B (n_2306), .C (n_4121), .D
       (\rs1_data[4]_39436 ), .Q (n_8494));
  AO22X2 g92821(.A (n_4147), .B (n_2258), .C (n_7686), .D (n_2303), .Q
       (n_8495));
  OA22X4 g92822(.A (n_4123), .B (n_2303), .C (n_2438), .D (n_2258), .Q
       (n_8496));
  AN21X1 g92823(.A (n_7684), .B (n_2303), .C (n_4188), .Q (n_8497));
  AO22X4 g92825(.A (n_8501), .B (n_2258), .C (n_7692), .D (n_2303), .Q
       (n_8499));
  NA3I2X4 g92827(.C (n_4024), .AN (n_8620), .BN (n_4008), .Q (n_8501));
  NO6I2X1 g92828(.C (n_3981), .D (n_3982), .E (n_3711), .F (n_3631),
       .AN (n_3729), .BN (n_3730), .Q (n_8502));
  NO6I2X4 g92830(.C (n_3917), .D (n_3911), .E (n_3563), .F (n_3540),
       .AN (n_3594), .BN (n_3595), .Q (n_8504));
  NO6I2X2 g92831(.C (n_3855), .D (n_3848), .E (n_3445), .F (n_3142),
       .AN (n_3460), .BN (n_3434), .Q (n_8505));
  NA3X2 g92832(.A (n_3611), .B (n_3612), .C (n_3912), .Q (n_8506));
  AN221X1 g92834(.A (n_3170), .B (n_7208), .C (n_3171), .D (n_7206), .E
       (n_3697), .Q (n_8508));
  NA3X1 g92835(.A (n_3476), .B (n_3486), .C (n_3857), .Q (n_8509));
  NA3X1 g92836(.A (n_3475), .B (n_3459), .C (n_3850), .Q (n_8510));
  NA3X2 g92837(.A (n_3421), .B (n_3410), .C (n_3841), .Q (n_8511));
  AN221X1 g92838(.A (n_3170), .B (n_6743), .C (n_3171), .D (n_6741), .E
       (n_3764), .Q (n_8512));
  AN221X1 g92839(.A (n_3170), .B (n_7146), .C (n_3171), .D (n_7144), .E
       (n_3763), .Q (n_8513));
  AN221X1 g92840(.A (n_3177), .B (n_6742), .C (n_3167), .D (n_6744), .E
       (n_3770), .Q (n_8514));
  AN221X1 g92841(.A (n_3175), .B (n_7143), .C (n_2300), .D (n_7141), .E
       (n_3750), .Q (n_8515));
  NA3I2X2 g92842(.C (n_8555), .AN (n_3248), .BN (n_3247), .Q (n_8516));
  AN221X1 g92843(.A (n_3159), .B (n_7027), .C (n_3161), .D (n_7025), .E
       (n_3583), .Q (n_8517));
  AN221X1 g92844(.A (n_3157), .B (n_6316), .C (n_3159), .D (n_6314), .E
       (n_3580), .Q (n_8518));
  AN221X1 g92845(.A (n_3159), .B (n_7213), .C (n_3161), .D (n_7211), .E
       (n_3576), .Q (n_8519));
  NA3I2X1 g92846(.C (n_8559), .AN (n_3274), .BN (n_2343), .Q (n_8520));
  AN211X1 g92848(.A (n_2587), .B (n_6473), .C (n_3525), .D (n_3232), .Q
       (n_8522));
  NO6I2X1 g92849(.C (n_2264), .D (n_8486), .E (n_8300), .F (n_2520),
       .AN (n_2592), .BN (n_8570), .Q (n_8523));
  OA21X2 g92852(.A (n_2530), .B (n_2590), .C (csr_data_out[21]), .Q
       (n_8526));
  OA21X2 g92853(.A (n_2546), .B (n_2590), .C (csr_data_out[20]), .Q
       (n_8527));
  OA21X2 g92854(.A (n_2532), .B (n_2590), .C (csr_data_out[18]), .Q
       (n_8528));
  AN221X1 g92855(.A (n_3057), .B (n_6913), .C (n_3064), .D (n_6912), .E
       (n_3488), .Q (n_8529));
  AN221X1 g92856(.A (n_3054), .B (n_6394), .C (n_3063), .D (n_6395), .E
       (n_3437), .Q (n_8530));
  AN221X1 g92857(.A (n_3104), .B (n_6328), .C (n_3055), .D (n_6325), .E
       (n_3413), .Q (n_8531));
  AN221X1 g92858(.A (n_3061), .B (n_7097), .C (n_2336), .D (n_7096), .E
       (n_3417), .Q (n_8532));
  AN221X1 g92859(.A (n_3105), .B (n_7198), .C (n_2339), .D (n_7197), .E
       (n_3510), .Q (n_8533));
  AN221X1 g92860(.A (n_3057), .B (n_6727), .C (n_3064), .D (n_6726), .E
       (n_3407), .Q (n_8534));
  AN221X1 g92861(.A (n_3054), .B (n_6828), .C (n_3063), .D (n_6829), .E
       (n_3277), .Q (n_8535));
  AN221X1 g92862(.A (n_3073), .B (n_7225), .C (n_3075), .D (n_7226), .E
       (n_3196), .Q (n_8536));
  AO222X2 g92863(.A (n_3073), .B (n_6636), .C (n_3075), .D (n_6637), .E
       (n_2339), .F (n_6639), .Q (n_8537));
  AN221X1 g92864(.A (n_3075), .B (n_6978), .C (n_2337), .D (n_6970), .E
       (n_3191), .Q (n_8538));
  AN222X1 g92865(.A (n_3073), .B (n_6543), .C (n_3075), .D (n_6544), .E
       (n_3051), .F (n_6548), .Q (n_8539));
  AN222X1 g92866(.A (n_3073), .B (n_6419), .C (n_3075), .D (n_6420), .E
       (n_3051), .F (n_6424), .Q (n_8540));
  AN221X1 g92867(.A (n_3073), .B (n_6884), .C (n_3075), .D (n_6885), .E
       (n_3210), .Q (n_8541));
  AO222X2 g92868(.A (n_3073), .B (n_7039), .C (n_3075), .D (n_7040), .E
       (n_3055), .F (n_7038), .Q (n_8542));
  AN22X1 g92869(.A (n_3177), .B (n_7114), .C (n_3175), .D (n_7112), .Q
       (n_8543));
  AO222X1 g92870(.A (n_3073), .B (n_6729), .C (n_3075), .D (n_6730), .E
       (n_3051), .F (n_6734), .Q (n_8544));
  AO222X2 g92871(.A (n_3073), .B (n_7132), .C (n_3075), .D (n_7133), .E
       (n_3051), .F (n_7137), .Q (n_8545));
  AN222X1 g92872(.A (n_3073), .B (n_7101), .C (n_3075), .D (n_7102), .E
       (n_3051), .F (n_7106), .Q (n_8546));
  AN222X1 g92873(.A (n_3073), .B (n_7008), .C (n_3075), .D (n_7009), .E
       (n_3052), .F (n_7013), .Q (n_8547));
  AO222X2 g92874(.A (n_3073), .B (n_7070), .C (n_3075), .D (n_7071), .E
       (n_3051), .F (n_7075), .Q (n_8548));
  AN221X1 g92876(.A (n_3054), .B (n_6487), .C (n_3063), .D (n_6488), .E
       (n_3251), .Q (n_8550));
  AN21X1 g92877(.A (n_3051), .B (n_6269), .C (n_3331), .Q (n_8551));
  AN21X1 g92878(.A (n_3175), .B (n_6678), .C (n_3259), .Q (n_8552));
  AN21X1 g92879(.A (n_3167), .B (n_6682), .C (n_3257), .Q (n_8553));
  AN21X1 g92880(.A (n_2587), .B (n_7000), .C (n_3314), .Q (n_8554));
  AN21X1 g92881(.A (n_2300), .B (n_6521), .C (n_3246), .Q (n_8555));
  AN22X1 g92882(.A (n_3156), .B (n_6534), .C (n_3154), .D (n_6532), .Q
       (n_8556));
  AN21X1 g92883(.A (n_3052), .B (n_6579), .C (n_3238), .Q (n_8557));
  AN22X1 g92884(.A (n_3157), .B (n_6657), .C (n_2587), .D (n_6659), .Q
       (n_8558));
  AN22X1 g92885(.A (n_3159), .B (n_7182), .C (n_2587), .D (n_7186), .Q
       (n_8559));
  AN22X1 g92886(.A (n_3107), .B (n_7157), .C (n_3066), .D (n_7156), .Q
       (n_8560));
  AN21X1 g92887(.A (n_3060), .B (n_6569), .C (n_3118), .Q (n_8561));
  AN21X1 g92889(.A (n_7282), .B (n_7303), .C (n_3040), .Q (n_8563));
  AO222X2 g92890(.A (n_2755), .B (csr_mcycle[1]), .C (n_2733), .D
       (csr_minstret[1]), .E (n_2727), .F (csr_mscratch[1]), .Q
       (n_8564));
  AO222X2 g92891(.A (n_2755), .B (csr_mcycle[3]), .C (n_2756), .D
       (csr_mcycle[35]), .E (n_2726), .F (csr_mtval[3]), .Q (n_8565));
  AO21X4 g92892(.A (n_8318), .B (n_2321), .C (n_2800), .Q (n_8566));
  AN22X1 g92893(.A (\rs1_data[3]_39426 ), .B (n_2589), .C (n_7680), .D
       (n_2311), .Q (n_8567));
  AN22X1 g92894(.A (\rs1_data[1]_39396 ), .B (n_2589), .C (n_7682), .D
       (n_2311), .Q (n_8568));
  AO21X1 g92895(.A (n_8054), .B (write_response), .C (n_2596), .Q
       (n_8569));
  NO3I1X4 g92896(.B (n_8482), .C (n_2491), .AN (n_2421), .Q (n_8570));
  AO21X4 g92897(.A (\rs1_data[24]_39336 ), .B (n_2589), .C (n_8525), .Q
       (n_8571));
  AN222X1 g92902(.A (n_7428), .B (n_159), .C (n_7518), .D (n_1101), .E
       (n_7519), .F (n_1100), .Q (n_8576));
  AN222X1 g92903(.A (n_7426), .B (n_159), .C (n_7514), .D (n_1101), .E
       (n_7515), .F (n_1100), .Q (n_8577));
  AN222X1 g92904(.A (n_7424), .B (n_159), .C (n_7510), .D (n_1101), .E
       (n_7511), .F (n_1100), .Q (n_8578));
  AN222X1 g92905(.A (n_7422), .B (n_159), .C (n_7506), .D (n_1101), .E
       (n_7507), .F (n_1100), .Q (n_8579));
  AND3X2 g92913(.A (n_2739), .B (n_2591), .C (n_1082), .Q (n_8587));
  NO3I2X4 g92914(.C (n_2509), .AN (n_1082), .BN (n_2739), .Q (n_8588));
  OA211X2 g92915(.A (n_781), .B (n_776), .C (n_533), .D (n_350), .Q
       (n_8589));
  OA211X1 g92917(.A (n_352), .B (alu_2nd_operand[1]), .C (n_691), .D
       (n_581), .Q (n_8591));
  NA3X1 g92918(.A (add_463_14_n_646), .B (add_463_14_n_760), .C
       (add_463_14_n_752), .Q (n_8592));
  OA221X2 g92919(.A (add_463_14_n_708), .B (add_463_14_n_840), .C
       (add_463_14_n_958), .D (add_463_14_n_948), .E
       (add_463_14_n_943), .Q (n_8593));
  AN21X1 g92920(.A (add_463_14_n_792), .B (add_463_14_n_780), .C
       (add_463_14_n_783), .Q (n_8594));
  AO221X2 g92921(.A (add_464_21_n_686), .B (add_464_21_n_749), .C
       (add_464_21_n_752), .D (add_464_21_n_944), .E
       (add_464_21_n_924), .Q (n_8595));
  NO3I2X1 g92922(.C (inc_ADD_UNS_OP_5_n_3583), .AN
       (inc_ADD_UNS_OP_5_n_3695), .BN (inc_ADD_UNS_OP_5_n_3697), .Q
       (n_8596));
  NA3X2 g92923(.A (inc_add_1345_58_1_n_3399), .B (csr_mcycle[2]), .C
       (csr_mcycle[3]), .Q (n_8597));
  NO3I1X2 g92924(.B (inc_add_1345_58_1_n_3455), .C
       (inc_ADD_UNS_OP5491_6_n_2657), .AN (inc_add_1345_58_1_n_3151),
       .Q (n_8598));
  NA3X2 g92925(.A (inc_add_1347_34_2_n_2561), .B (csr_mcycle[2]), .C
       (csr_mcycle[3]), .Q (n_8599));
  AND6X2 g92926(.A (inc_ADD_UNS_OP5492_3_n_2504), .B
       (inc_ADD_UNS_OP5492_3_n_2574), .C (csr_minstret[22]), .D
       (csr_minstret[23]), .E (csr_minstret[25]), .F
       (csr_minstret[24]), .Q (n_8600));
  AND4X2 g92928(.A (n_5871), .B (n_8671), .C (n_8429), .D (n_5884), .Q
       (n_8602));
  NO6I4X1 g92929(.E (n_5486), .F (n_5484), .AN (n_5529), .BN (n_5539),
       .CN (n_5847), .DN (n_5841), .Q (n_8603));
  AND5X1 g92930(.A (n_5419), .B (n_5541), .C (n_4822), .D (n_4821), .E
       (n_5528), .Q (n_8604));
  OR4X2 g92931(.A (n_5731), .B (n_5723), .C (n_5667), .D (n_5714), .Q
       (n_8605));
  NA5I2X2 g92932(.C (n_5519), .D (n_5513), .E (n_8458), .AN (n_5160),
       .BN (n_5161), .Q (n_8606));
  OR4X1 g92933(.A (n_4848), .B (n_5641), .C (n_5559), .D (n_5553), .Q
       (n_8607));
  OR4X1 g92934(.A (n_5468), .B (n_5481), .C (n_5469), .D (n_5480), .Q
       (n_8608));
  NA5I1X4 g92935(.B (n_5072), .C (n_5079), .D (n_5438), .E (n_5446),
       .AN (n_5454), .Q (n_8609));
  AND4X1 g92936(.A (n_5389), .B (n_5390), .C (n_5393), .D (n_5394), .Q
       (n_8610));
  NO6I2X4 g92937(.C (n_4841), .D (n_4842), .E (n_4835), .F (n_4836),
       .AN (n_5372), .BN (n_5359), .Q (n_8611));
  AND4X1 g92938(.A (n_5362), .B (n_5352), .C (n_8476), .D (n_5351), .Q
       (n_8612));
  AND4X1 g92939(.A (n_5353), .B (n_5354), .C (n_8475), .D (n_8474), .Q
       (n_8613));
  AND4X2 g92941(.A (n_5330), .B (n_5331), .C (n_5320), .D (n_5321), .Q
       (n_8615));
  AND4X2 g92942(.A (n_5183), .B (n_5177), .C (n_5156), .D (n_5157), .Q
       (n_8616));
  AN221X1 g92943(.A (n_4452), .B (n_6623), .C (n_4883), .D (n_6624), .E
       (n_5456), .Q (n_8617));
  AN22X1 g92944(.A (n_4884), .B (n_6639), .C (n_4889), .D (n_6638), .Q
       (n_8618));
  OR4X2 g92945(.A (n_3996), .B (n_3956), .C (n_4058), .D (n_4030), .Q
       (n_8619));
  OR4X2 g92946(.A (n_3557), .B (n_3544), .C (n_3543), .D (n_3554), .Q
       (n_8620));
  OR4X2 g92947(.A (n_3236), .B (n_3117), .C (n_3254), .D (n_3241), .Q
       (n_8621));
  AO22X4 g92948(.A (n_2655), .B (csr_data_out[16]), .C (n_6132), .D
       (n_2589), .Q (n_8622));
  OR4X1 g92949(.A (n_325), .B (n_324), .C (n_327), .D (n_326), .Q
       (n_8623));
  NO6I2X4 g92950(.C (n_4843), .D (n_5635), .E (n_8456), .F (n_5650),
       .AN (n_8434), .BN (n_5848), .Q (n_8624));
  NO5I3X2 g92951(.D (n_4773), .E (n_4774), .AN (n_5336), .BN (n_5337),
       .CN (n_5417), .Q (n_8625));
  ON21X1 g92978(.A (n_8652), .B (n_4137), .C (n_4229), .Q (n_8653));
  NO2X1 g92979(.A (n_2379), .B (n_6135), .Q (n_8652));
  OA21X4 g92980(.A (n_2432), .B (n_2588), .C (n_8654), .Q (n_8655));
  ON21X1 g92981(.A (n_2542), .B (n_2590), .C (csr_data_out[23]), .Q
       (n_8654));
  OA21X2 g92982(.A (n_2429), .B (n_2588), .C (n_8656), .Q (n_8657));
  ON21X1 g92983(.A (n_2536), .B (n_2590), .C (csr_data_out[11]), .Q
       (n_8656));
  NA2X4 g92984(.A (n_8658), .B (n_2621), .Q (n_8659));
  ON21X1 g92985(.A (n_2478), .B (instruction[22]), .C
       (instruction[23]), .Q (n_8658));
  NA2X2 g92986(.A (n_8660), .B (n_175), .Q (n_8661));
  EO2X1 g92987(.A (inc_add_1343_59_4_n_3423), .B (csr_mcycle[63]), .Q
       (n_8660));
  NA3I1X2 g92988(.B (n_8450), .C (n_8662), .AN (n_5108), .Q (n_8663));
  AN21X1 g92989(.A (n_4741), .B (n_6598), .C (n_5107), .Q (n_8662));
  HAX2 g92990(.A (csr_mcause_code[0]), .B (csr_mtvec[2]), .S (n_8664),
       .CO (n_8665));
  DFRQX2 prev_write_request_reg(.C (rc_gclk), .D (n_1490), .Q (n_8054));
  DFRQX1 \program_counter_reg[0] (.C (rc_gclk_199879), .D (n_1486), .Q
       (program_counter[0]));
  DFRQX1 csr_mstatus_mie_reg(.C (rc_gclk), .D (n_2057), .Q (n_7275));
  DFRQX1 \program_counter_reg[2] (.C (rc_gclk_199879), .D (n_1464), .Q
       (program_counter[2]));
  DFRQX1 \program_counter_reg[3] (.C (rc_gclk_199879), .D (n_1461), .Q
       (program_counter[3]));
  DFRQX1 \program_counter_reg[4] (.C (rc_gclk_199879), .D (n_1460), .Q
       (program_counter[4]));
  DFRQX1 \program_counter_reg[5] (.C (rc_gclk_199879), .D (n_1459), .Q
       (program_counter[5]));
  DFRQX1 \program_counter_reg[7] (.C (rc_gclk_199879), .D (n_1457), .Q
       (program_counter[7]));
  DFRQX1 \program_counter_reg[6] (.C (rc_gclk_199879), .D (n_1458), .Q
       (program_counter[6]));
  DFRQX1 \program_counter_reg[8] (.C (rc_gclk_199879), .D (n_1456), .Q
       (program_counter[8]));
  DFRQX1 \program_counter_reg[9] (.C (rc_gclk_199879), .D (n_1455), .Q
       (program_counter[9]));
  DFRQX1 \program_counter_reg[11] (.C (rc_gclk_199879), .D (n_1484), .Q
       (program_counter[11]));
  DFRQX1 \program_counter_reg[10] (.C (rc_gclk_199879), .D (n_1485), .Q
       (program_counter[10]));
  DFRQX1 \program_counter_reg[12] (.C (rc_gclk_199879), .D (n_1483), .Q
       (program_counter[12]));
  DFRQX1 \program_counter_reg[13] (.C (rc_gclk_199879), .D (n_1482), .Q
       (program_counter[13]));
  DFRQX1 \program_counter_reg[15] (.C (rc_gclk_199879), .D (n_1480), .Q
       (program_counter[15]));
  DFRQX1 \program_counter_reg[14] (.C (rc_gclk_199879), .D (n_1481), .Q
       (program_counter[14]));
  DFRQX1 \program_counter_reg[16] (.C (rc_gclk_199879), .D (n_1479), .Q
       (program_counter[16]));
  DFRQX1 \program_counter_reg[17] (.C (rc_gclk_199879), .D (n_1478), .Q
       (program_counter[17]));
  DFRQX1 \program_counter_reg[19] (.C (rc_gclk_199879), .D (n_1476), .Q
       (program_counter[19]));
  DFRQX1 \program_counter_reg[18] (.C (rc_gclk_199879), .D (n_1477), .Q
       (program_counter[18]));
  DFRQX1 \program_counter_reg[20] (.C (rc_gclk_199879), .D (n_1474), .Q
       (program_counter[20]));
  DFRQX1 \program_counter_reg[21] (.C (rc_gclk_199879), .D (n_1473), .Q
       (program_counter[21]));
  DFRQX1 \program_counter_reg[23] (.C (rc_gclk_199879), .D (n_1471), .Q
       (program_counter[23]));
  DFRQX1 \program_counter_reg[22] (.C (rc_gclk_199879), .D (n_1472), .Q
       (program_counter[22]));
  DFRQX1 \program_counter_reg[24] (.C (rc_gclk_199879), .D (n_1470), .Q
       (program_counter[24]));
  DFRQX1 \program_counter_reg[25] (.C (rc_gclk_199879), .D (n_1469), .Q
       (program_counter[25]));
  DFRQX1 \program_counter_reg[27] (.C (rc_gclk_199879), .D (n_1467), .Q
       (program_counter[27]));
  DFRQX1 \program_counter_reg[26] (.C (rc_gclk_199879), .D (n_1468), .Q
       (program_counter[26]));
  DFRQX1 \program_counter_reg[28] (.C (rc_gclk_199879), .D (n_1466), .Q
       (program_counter[28]));
  DFRQX1 \program_counter_reg[29] (.C (rc_gclk_199879), .D (n_1465), .Q
       (program_counter[29]));
  DFRQX1 \program_counter_reg[30] (.C (rc_gclk_199879), .D (n_1463), .Q
       (program_counter[30]));
  DFRQX1 \program_counter_reg[31] (.C (rc_gclk_199879), .D (n_1462), .Q
       (program_counter[31]));
  DFRQX1 \csr_mcause_code_reg[4] (.C (rc_gclk_199992), .D (n_7304), .Q
       (csr_mcause_code[4]));
  DFRQX1 \csr_mcause_code_reg[3] (.C (rc_gclk_199992), .D (n_2256), .Q
       (csr_mcause_code[3]));
  DFRQX1 \csr_mcause_code_reg[1] (.C (rc_gclk_199992), .D (n_2254), .Q
       (csr_mcause_code[1]));
  DFRQX1 \csr_mcause_code_reg[0] (.C (rc_gclk_199992), .D (n_2257), .Q
       (csr_mcause_code[0]));
  DFRQX1 \csr_mcycle_reg[32] (.C (clock), .D (n_2202), .Q
       (csr_mcycle[32]));
  DFRQX1 \csr_minstret_reg[32] (.C (rc_gclk), .D (n_2102), .Q
       (csr_minstret[32]));
  DFRQX1 \csr_mcycle_reg[42] (.C (clock), .D (n_2191), .Q
       (csr_mcycle[42]));
  DFRQX1 \csr_minstret_reg[42] (.C (rc_gclk), .D (n_2091), .Q
       (csr_minstret[42]));
  DFRQX1 \csr_mcycle_reg[10] (.C (clock), .D (n_2226), .Q
       (csr_mcycle[10]));
  DFRQX1 \csr_minstret_reg[10] (.C (rc_gclk), .D (n_2126), .Q
       (csr_minstret[10]));
  DFRQX1 \csr_mcycle_reg[43] (.C (clock), .D (n_2190), .Q
       (csr_mcycle[43]));
  DFRQX1 \csr_minstret_reg[43] (.C (rc_gclk), .D (n_2090), .Q
       (csr_minstret[43]));
  DFRQX1 \csr_mcycle_reg[44] (.C (clock), .D (n_2189), .Q
       (csr_mcycle[44]));
  DFRQX1 \csr_minstret_reg[44] (.C (rc_gclk), .D (n_2089), .Q
       (csr_minstret[44]));
  DFRQX1 \csr_mcycle_reg[45] (.C (clock), .D (n_2188), .Q
       (csr_mcycle[45]));
  DFRQX1 \csr_minstret_reg[45] (.C (rc_gclk), .D (n_2088), .Q
       (csr_minstret[45]));
  DFRQX1 \csr_mcycle_reg[46] (.C (clock), .D (n_2187), .Q
       (csr_mcycle[46]));
  DFRQX1 \csr_minstret_reg[46] (.C (rc_gclk), .D (n_2087), .Q
       (csr_minstret[46]));
  DFRQX1 \csr_mcycle_reg[47] (.C (clock), .D (n_2186), .Q
       (csr_mcycle[47]));
  DFRQX1 \csr_minstret_reg[47] (.C (rc_gclk), .D (n_2086), .Q
       (csr_minstret[47]));
  DFRQX1 \csr_minstret_reg[48] (.C (rc_gclk), .D (n_2085), .Q
       (csr_minstret[48]));
  DFRQX1 \csr_mcycle_reg[16] (.C (clock), .D (n_2220), .Q
       (csr_mcycle[16]));
  DFRQX1 \csr_minstret_reg[16] (.C (rc_gclk), .D (n_2120), .Q
       (csr_minstret[16]));
  DFRQX1 \csr_mcycle_reg[49] (.C (clock), .D (n_2184), .Q
       (csr_mcycle[49]));
  DFRQX1 \csr_mcycle_reg[17] (.C (clock), .D (n_2219), .Q
       (csr_mcycle[17]));
  DFRQX1 \csr_minstret_reg[17] (.C (rc_gclk), .D (n_2119), .Q
       (csr_minstret[17]));
  DFRQX1 \csr_mcycle_reg[18] (.C (clock), .D (n_2218), .Q
       (csr_mcycle[18]));
  DFRQX1 \csr_minstret_reg[18] (.C (rc_gclk), .D (n_2118), .Q
       (csr_minstret[18]));
  DFRQX1 \csr_mcycle_reg[51] (.C (clock), .D (n_2181), .Q
       (csr_mcycle[51]));
  DFRQX1 \csr_mcycle_reg[33] (.C (clock), .D (n_2201), .Q
       (csr_mcycle[33]));
  DFRQX1 \csr_mcycle_reg[52] (.C (clock), .D (n_2180), .Q
       (csr_mcycle[52]));
  DFRQX1 \csr_mcycle_reg[20] (.C (clock), .D (n_2215), .Q
       (csr_mcycle[20]));
  DFRQX1 \csr_minstret_reg[20] (.C (rc_gclk), .D (n_2115), .Q
       (csr_minstret[20]));
  DFRQX1 \csr_minstret_reg[53] (.C (rc_gclk), .D (n_2079), .Q
       (csr_minstret[53]));
  DFRQX1 \csr_mcycle_reg[55] (.C (clock), .D (n_2177), .Q
       (csr_mcycle[55]));
  DFRQX1 \csr_minstret_reg[55] (.C (rc_gclk), .D (n_2077), .Q
       (csr_minstret[55]));
  DFRQX1 \csr_mcycle_reg[57] (.C (clock), .D (n_2175), .Q
       (csr_mcycle[57]));
  DFRQX1 \csr_minstret_reg[57] (.C (rc_gclk), .D (n_2075), .Q
       (csr_minstret[57]));
  DFRQX1 \csr_mcycle_reg[59] (.C (clock), .D (n_2173), .Q
       (csr_mcycle[59]));
  DFRQX1 \csr_minstret_reg[59] (.C (rc_gclk), .D (n_2073), .Q
       (csr_minstret[59]));
  DFRQX1 \csr_mcycle_reg[34] (.C (clock), .D (n_2200), .Q
       (csr_mcycle[34]));
  DFRQX1 \csr_minstret_reg[34] (.C (rc_gclk), .D (n_2100), .Q
       (csr_minstret[34]));
  DFRQX1 \csr_minstret_reg[2] (.C (rc_gclk), .D (n_2105), .Q
       (csr_minstret[2]));
  DFRQX1 \csr_mcycle_reg[30] (.C (clock), .D (n_2204), .Q
       (csr_mcycle[30]));
  DFRQX1 \csr_mcycle_reg[62] (.C (clock), .D (n_2169), .Q
       (csr_mcycle[62]));
  DFRSQX1 \csr_mcycle_reg[35] (.SN (1'b1), .C (clock), .D (n_2199), .Q
       (csr_mcycle[35]));
  DFRQX1 \csr_minstret_reg[36] (.C (rc_gclk), .D (n_2098), .Q
       (csr_minstret[36]));
  DFRQX1 \csr_minstret_reg[37] (.C (rc_gclk), .D (n_2097), .Q
       (csr_minstret[37]));
  DFRQX1 \csr_mcycle_reg[38] (.C (clock), .D (n_2196), .Q
       (csr_mcycle[38]));
  DFRQX1 \csr_minstret_reg[38] (.C (rc_gclk), .D (n_2096), .Q
       (csr_minstret[38]));
  DFRQX1 \csr_mcycle_reg[6] (.C (clock), .D (n_2167), .Q
       (csr_mcycle[6]));
  DFRQX1 \csr_mcycle_reg[39] (.C (clock), .D (n_2195), .Q
       (csr_mcycle[39]));
  DFRQX1 \csr_minstret_reg[39] (.C (rc_gclk), .D (n_2095), .Q
       (csr_minstret[39]));
  DFRQX1 \csr_mcycle_reg[40] (.C (clock), .D (n_2193), .Q
       (csr_mcycle[40]));
  DFRQX1 \csr_minstret_reg[40] (.C (rc_gclk), .D (n_2093), .Q
       (csr_minstret[40]));
  DFRQX1 \csr_mcycle_reg[8] (.C (clock), .D (n_2165), .Q
       (csr_mcycle[8]));
  DFRQX1 \csr_minstret_reg[8] (.C (rc_gclk), .D (n_2065), .Q
       (csr_minstret[8]));
  DFRQX1 \csr_mcycle_reg[41] (.C (clock), .D (n_2192), .Q
       (csr_mcycle[41]));
  DFRQX1 \csr_minstret_reg[41] (.C (rc_gclk), .D (n_2092), .Q
       (csr_minstret[41]));
  DFRQX1 \csr_minstret_reg[9] (.C (rc_gclk), .D (n_2064), .Q
       (csr_minstret[9]));
  INX2 g93180(.A (n_2939), .Q (n_2940));
  AND2X2 g93182(.A (n_5434), .B (n_5447), .Q (n_5807));
  INX2 g93184(.A (n_4489), .Q (n_4750));
  INX2 g93186(.A (n_2314), .Q (n_2614));
  AND2X1 g93190(.A (n_4723), .B (n_8485), .Q (n_8257));
  AND6X1 g93194(.A (n_8413), .B (n_5903), .C (n_5717), .D (n_5725), .E
       (n_5704), .F (n_5696), .Q (n_6073));
  AND6X1 g93196(.A (n_8414), .B (n_5904), .C (n_5718), .D (n_5726), .E
       (n_5705), .F (n_5697), .Q (n_6072));
  NO5X2 g93198(.A (n_5784), .B (n_4991), .C (n_4992), .D (n_4993), .E
       (n_4994), .Q (n_8398));
  AO321X1 add_464_21_g93200(.A (add_464_21_n_941), .B
       (add_464_21_n_708), .C (add_464_21_n_637), .D
       (add_464_21_n_941), .E (add_464_21_n_686), .F
       (add_464_21_n_930), .Q (add_464_21_n_605));
  AO321X1 add_464_21_g93202(.A (add_464_21_n_946), .B
       (add_464_21_n_730), .C (add_464_21_n_637), .D
       (add_464_21_n_946), .E (add_464_21_n_701), .F
       (add_464_21_n_919), .Q (add_464_21_n_611));
  ON21X2 g93204(.A (n_3044), .B (n_4115), .C (n_4293), .Q
       (write_data[31]));
  ON21X2 g93206(.A (n_3044), .B (n_4114), .C (n_4292), .Q
       (write_data[30]));
  ON21X2 g93208(.A (n_3044), .B (n_4131), .C (n_4291), .Q
       (write_data[29]));
  ON21X2 g93210(.A (n_3044), .B (n_4121), .C (n_4290), .Q
       (write_data[28]));
  ON21X2 g93212(.A (n_3044), .B (n_2365), .C (n_4289), .Q
       (write_data[27]));
  ON21X2 g93214(.A (n_3044), .B (n_4123), .C (n_4288), .Q
       (write_data[26]));
  ON21X2 g93216(.A (n_3044), .B (n_2366), .C (n_4287), .Q
       (write_data[25]));
  ON21X2 g93218(.A (n_3044), .B (n_4116), .C (n_4286), .Q
       (write_data[24]));
  AND2X1 add_463_14_g93220(.A (add_463_14_n_759), .B
       (add_463_14_n_762), .Q (add_463_14_n_726));
  INX2 g93222(.A (n_8054), .Q (n_4526));
  AND2X2 g93224(.A (n_7825), .B (n_2721), .Q (n_2800));
  ON21X1 g93226(.A (n_5230), .B (n_4470), .C (n_5228), .Q (n_7687));
  OA21X1 g93228(.A (n_2534), .B (n_2590), .C (csr_data_out[24]), .Q
       (n_8525));
  OA221X1 g93230(.A (n_734), .B (n_8591), .C (n_378), .D (n_340), .E
       (n_635), .Q (n_357));
  AND2X2 g93232(.A (take_trap_39229), .B (n_7861), .Q (n_158));
  INX2 g93234(.A (n_4687), .Q (n_4688));
  INX2 g93236(.A (n_4648), .Q (n_4649));
  INX2 g93238(.A (n_2304), .Q (n_2305));
  NO2I1X2 g93240(.B (n_2490), .AN (n_2431), .Q (n_2521));
  NO2X4 g93241(.A (n_7862), .B (n_8297), .Q (n_8666));
  AN221X1 g93244(.A (n_4888), .B (n_7196), .C (n_4884), .D (n_7197), .E
       (n_5710), .Q (n_8669));
  AN221X1 g93245(.A (n_4884), .B (n_7104), .C (n_4888), .D (n_7103), .E
       (n_5627), .Q (n_8670));
  AN221X1 g93246(.A (n_4870), .B (n_7160), .C (n_4868), .D (n_7159), .E
       (n_5492), .Q (n_8671));
  AO22X2 g93248(.A (n_4500), .B (n_7181), .C (n_4883), .D (n_7182), .Q
       (n_8673));
  AO22X2 g93249(.A (n_4878), .B (n_6456), .C (n_4506), .D (n_6457), .Q
       (n_8674));
  AO22X2 g93250(.A (n_4484), .B (n_6501), .C (n_4744), .D (n_6502), .Q
       (n_8675));
  AO22X2 g93251(.A (n_4465), .B (prev_instruction[12]), .C (n_4467), .D
       (read_data[12]), .Q (n_8676));
  AO22X4 g93252(.A (n_2367), .B (n_2258), .C (n_2437), .D (n_2303), .Q
       (n_8677));
  AN221X1 g93253(.A (n_3170), .B (n_7053), .C (n_3171), .D (n_7051), .E
       (n_3755), .Q (n_8678));
  AN221X1 g93255(.A (n_3075), .B (n_6513), .C (n_3073), .D (n_6512), .E
       (n_3134), .Q (n_8680));
  AN221X1 g93256(.A (n_3073), .B (n_6853), .C (n_3075), .D (n_6854), .E
       (n_3133), .Q (n_8681));
  AN21X1 g93257(.A (n_3052), .B (n_6455), .C (n_3237), .Q (n_8682));
  AN222X1 g93262(.A (n_7421), .B (n_159), .C (n_7504), .D (n_1101), .E
       (n_7505), .F (n_1100), .Q (n_8687));
  AN222X1 g93263(.A (n_7419), .B (n_159), .C (n_7500), .D (n_1101), .E
       (n_7501), .F (n_1100), .Q (n_8688));
  AN222X1 g93264(.A (n_7417), .B (n_159), .C (n_7496), .D (n_1101), .E
       (n_7497), .F (n_1100), .Q (n_8689));
  AN222X1 g93265(.A (n_7415), .B (n_159), .C (n_7492), .D (n_1101), .E
       (n_7493), .F (n_1100), .Q (n_8690));
  AN222X1 g93266(.A (n_7410), .B (n_159), .C (n_7482), .D (n_1101), .E
       (n_7483), .F (n_1100), .Q (n_8691));
  AN222X1 g93267(.A (n_7409), .B (n_159), .C (n_7480), .D (n_1101), .E
       (n_7481), .F (n_1100), .Q (n_8692));
  AND4X1 g93269(.A (n_5503), .B (n_5488), .C (n_5347), .D (n_5510), .Q
       (n_8694));
  OR4X2 g93270(.A (n_5482), .B (n_4788), .C (n_8462), .D (n_8461), .Q
       (n_8695));
  AN222X1 g93271(.A (n_4741), .B (n_6319), .C (n_4903), .D (n_6324), .E
       (n_4861), .F (n_6320), .Q (n_8696));
  AND4X2 g93272(.A (n_5182), .B (n_5176), .C (n_5154), .D (n_5155), .Q
       (n_8697));
  OR4X2 g93273(.A (n_5090), .B (n_5091), .C (n_5070), .D (n_5086), .Q
       (n_8698));
  OR4X2 g93274(.A (n_4817), .B (n_4818), .C (n_4815), .D (n_4816), .Q
       (n_8699));
  OR4X2 g93275(.A (n_3941), .B (n_3936), .C (n_3942), .D (n_8520), .Q
       (n_8700));
  AN222X1 g93276(.A (n_3051), .B (n_6300), .C (n_3073), .D (n_6295), .E
       (n_3075), .F (n_6296), .Q (n_8701));
  AN211X1 g93277(.A (n_4741), .B (n_6505), .C (n_5106), .D (n_5102), .Q
       (n_8702));
  DFRQX2 prev_load_request_reg(.C (rc_gclk), .D (n_1554), .Q
       (prev_load_request));
  DFRQX1 \csr_mcause_code_reg[2] (.C (rc_gclk_199992), .D (n_2252), .Q
       (csr_mcause_code[2]));
  DFRQX1 \csr_mcycle_reg[37] (.C (clock), .D (n_2197), .Q
       (csr_mcycle[37]));
  AND2X1 g93298(.A (n_4723), .B (n_8486), .Q (n_8258));
endmodule

